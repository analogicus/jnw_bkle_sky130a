magic
tech sky130A
magscale 1 1
timestamp 1746183817
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 5765 5358 5815
<< locali >>
rect -100 -100 5358 -50
<< m1 >>
rect -100 -50 -50 5765
<< m1 >>
rect 5308 -50 5358 5765
<< locali >>
rect -107 5758 -43 5822
<< m1 >>
rect -107 5758 -43 5822
<< viali >>
rect -100 5765 -50 5815
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 5301 5758 5365 5822
<< m1 >>
rect 5301 5758 5365 5822
<< viali >>
rect 5308 5765 5358 5815
<< locali >>
rect 5301 -107 5365 -43
<< m1 >>
rect 5301 -107 5365 -43
<< viali >>
rect 5308 -100 5358 -50
<< locali >>
rect -200 5865 5458 5915
<< locali >>
rect -200 -200 5458 -150
<< m1 >>
rect -200 -150 -150 5865
<< m1 >>
rect 5408 -150 5458 5865
<< locali >>
rect -207 5858 -143 5922
<< m1 >>
rect -207 5858 -143 5922
<< viali >>
rect -200 5865 -150 5915
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 5401 5858 5465 5922
<< m1 >>
rect 5401 5858 5465 5922
<< viali >>
rect 5408 5865 5458 5915
<< locali >>
rect 5401 -207 5465 -143
<< m1 >>
rect 5401 -207 5465 -143
<< viali >>
rect 5408 -200 5458 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 5308 5765
<< labels >>
flabel locali s -100 5765 5358 5815 0 FreeSans 400 0 0 0 VDD
port 57 nsew signal bidirectional
flabel locali s -200 5865 5458 5915 0 FreeSans 400 0 0 0 VSS
port 58 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744372385
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1400
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1160
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 1400
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 1160
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1296 0 1 1800
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1296 0 1 2200
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1800
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 2200
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1296 0 1 1400
box 0 0 832 400
use JNWATR_PCH_12C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1400
box 0 0 832 400
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 600
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1000
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT mirror2_MN4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 360
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 600
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 1000
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT mirror2_MN3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 360
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 2200
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 1800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3280 0 1 2200
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1296 0 1 1000
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1296 0 1 760
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1000
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 760
box 0 0 832 240
<< locali >>
rect 150 2550 4106 2650
<< locali >>
rect 150 150 4106 250
<< m1 >>
rect 150 250 250 2550
<< m1 >>
rect 4006 250 4106 2550
<< locali >>
rect 143 2543 257 2657
<< m1 >>
rect 143 2543 257 2657
<< viali >>
rect 150 2550 250 2650
<< locali >>
rect 143 143 257 257
<< m1 >>
rect 143 143 257 257
<< viali >>
rect 150 150 250 250
<< locali >>
rect 3999 2543 4113 2657
<< m1 >>
rect 3999 2543 4113 2657
<< viali >>
rect 4006 2550 4106 2650
<< locali >>
rect 3999 143 4113 257
<< m1 >>
rect 3999 143 4113 257
<< viali >>
rect 4006 150 4106 250
<< locali >>
rect 0 2700 4256 2800
<< locali >>
rect 0 0 4256 100
<< m1 >>
rect 0 100 100 2700
<< m1 >>
rect 4156 100 4256 2700
<< locali >>
rect -7 2693 107 2807
<< m1 >>
rect -7 2693 107 2807
<< viali >>
rect 0 2700 100 2800
<< locali >>
rect -7 -7 107 107
<< m1 >>
rect -7 -7 107 107
<< viali >>
rect 0 0 100 100
<< locali >>
rect 4149 2693 4263 2807
<< m1 >>
rect 4149 2693 4263 2807
<< viali >>
rect 4156 2700 4256 2800
<< locali >>
rect 4149 -7 4263 107
<< m1 >>
rect 4149 -7 4263 107
<< viali >>
rect 4156 0 4256 100
<< locali >>
rect 1248 2100 1536 2140
<< locali >>
rect 1888 1980 2048 2020
<< locali >>
rect 2080 2100 2368 2140
<< locali >>
rect 1248 1700 1536 1740
<< locali >>
rect 2080 1700 2368 1740
<< locali >>
rect 2720 1580 2880 1620
<< locali >>
rect 352 900 640 940
<< locali >>
rect 3232 900 3520 940
<< locali >>
rect 3616 780 3776 820
<< locali >>
rect 352 2100 640 2140
<< locali >>
rect 736 1980 896 2020
<< locali >>
rect 3232 2100 3520 2140
<< locali >>
rect 1248 1300 1536 1340
<< locali >>
rect 2080 1300 2368 1340
<< locali >>
rect 150 2272 4106 2368
<< locali >>
rect 143 2265 257 2375
<< m1 >>
rect 143 2265 257 2375
<< viali >>
rect 150 2272 250 2368
<< locali >>
rect 3999 2265 4113 2375
<< m1 >>
rect 3999 2265 4113 2375
<< viali >>
rect 4006 2272 4106 2368
<< locali >>
rect 0 432 4256 528
<< locali >>
rect -7 425 107 535
<< m1 >>
rect -7 425 107 535
<< viali >>
rect 0 432 100 528
<< locali >>
rect 4149 425 4263 535
<< m1 >>
rect 4149 425 4263 535
<< viali >>
rect 4156 432 4256 528
<< labels >>
flabel locali s 0 2700 4256 2800 0 FreeSans 400 0 0 0 VSS
port 5 nsew signal bidirectional
flabel locali s 150 2550 4106 2650 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 2
timestamp 1744122265
<< metal4 >>
rect -849 539 849 580
rect -849 -539 593 539
rect 829 -539 849 539
rect -849 -580 849 -539
<< via4 >>
rect 593 -539 829 539
<< mimcap2 >>
rect -769 460 231 500
rect -769 -460 -729 460
rect 191 -460 231 460
rect -769 -500 231 -460
<< mimcap2contact >>
rect -729 -460 191 460
<< metal5 >>
rect -753 -460 -729 460
rect 191 -460 215 460
rect -753 -484 215 -460
rect 551 -539 593 539
rect 829 -539 871 539
rect 551 -581 871 -539
<< labels >>
flabel metal5 s -849 -539 539 100 0 FreeSans 800 0 0 0 A
port 1 nsew signal bidirectional
flabel metal4 s 0 0 680 100 0 FreeSans 800 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2000 2000
<< end >>

magic
tech sky130A
magscale 1 1
timestamp 1748204603
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 4158 7706 4208
<< locali >>
rect -100 -100 7706 -50
<< m1 >>
rect -100 -50 -50 4158
<< m1 >>
rect 7656 -50 7706 4158
<< locali >>
rect -107 4151 -43 4215
<< m1 >>
rect -107 4151 -43 4215
<< viali >>
rect -100 4158 -50 4208
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 7649 4151 7713 4215
<< m1 >>
rect 7649 4151 7713 4215
<< viali >>
rect 7656 4158 7706 4208
<< locali >>
rect 7649 -107 7713 -43
<< m1 >>
rect 7649 -107 7713 -43
<< viali >>
rect 7656 -100 7706 -50
<< locali >>
rect -200 4258 7806 4308
<< locali >>
rect -200 -200 7806 -150
<< m1 >>
rect -200 -150 -150 4258
<< m1 >>
rect 7756 -150 7806 4258
<< locali >>
rect -207 4251 -143 4315
<< m1 >>
rect -207 4251 -143 4315
<< viali >>
rect -200 4258 -150 4308
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 7749 4251 7813 4315
<< m1 >>
rect 7749 4251 7813 4315
<< viali >>
rect 7756 4258 7806 4308
<< locali >>
rect 7749 -207 7813 -143
<< m1 >>
rect 7749 -207 7813 -143
<< viali >>
rect 7756 -200 7806 -150
use COMP4 U2_COMP4 
transform 1 0 0 0 1 0
box 0 0 2298 4158
<< labels >>
flabel locali s -200 4258 7806 4308 0 FreeSans 400 0 0 0 VDD
port 191 nsew signal bidirectional
flabel locali s -100 4158 7706 4208 0 FreeSans 400 0 0 0 VSS
port 192 nsew signal bidirectional
<< properties >>
<< end >>
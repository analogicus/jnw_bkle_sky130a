magic
tech sky130A
magscale 1 1
timestamp 1746029693
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 1700
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 1460
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 1700
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 1460
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 2100
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 2100
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 2900
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 2900
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 2500
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 2500
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 3300
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 3700
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 3300
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 3700
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 500
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 900
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 260
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 500
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 900
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 260
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2320
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4170
box 0 0 2236 1720
<< m1 >>
rect 3009 1873 3055 1927
<< m2 >>
rect 3009 1873 3055 1927
<< via1 >>
rect 3016 1880 3048 1920
<< m1 >>
rect 3585 1873 3631 1927
<< m2 >>
rect 3585 1873 3631 1927
<< via1 >>
rect 3592 1880 3624 1920
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< m3 >>
rect 3585 2273 3631 2327
<< via2 >>
rect 3592 2280 3624 2320
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< via1 >>
rect 3016 2280 3048 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< m3 >>
rect 3009 2273 3055 2327
<< via2 >>
rect 3016 2280 3048 2320
<< via1 >>
rect 3016 2280 3048 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< via1 >>
rect 3016 2280 3048 2320
<< m1 >>
rect 3585 3073 3631 3127
<< m2 >>
rect 3585 3073 3631 3127
<< via1 >>
rect 3592 3080 3624 3120
<< m1 >>
rect 3009 3073 3055 3127
<< m2 >>
rect 3009 3073 3055 3127
<< via1 >>
rect 3016 3080 3048 3120
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< m3 >>
rect 3009 2673 3055 2727
<< via2 >>
rect 3016 2680 3048 2720
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< via1 >>
rect 3592 2680 3624 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< m3 >>
rect 3585 2673 3631 2727
<< via2 >>
rect 3592 2680 3624 2720
<< via1 >>
rect 3592 2680 3624 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< via1 >>
rect 3592 2680 3624 2720
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< m3 >>
rect 3841 2913 3951 2967
<< via2 >>
rect 3848 2920 3944 2960
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< m3 >>
rect 3841 2913 3951 2967
<< via2 >>
rect 3848 2920 3944 2960
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< m3 >>
rect 3265 2913 3375 2967
<< via2 >>
rect 3272 2920 3368 2960
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< m3 >>
rect 3265 2913 3375 2967
<< via2 >>
rect 3272 2920 3368 2960
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< m3 >>
rect 3265 2513 3375 2567
<< via2 >>
rect 3272 2520 3368 2560
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< m3 >>
rect 3265 2513 3375 2567
<< via2 >>
rect 3272 2520 3368 2560
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3841 2513 3951 2567
<< m2 >>
rect 3841 2513 3951 2567
<< m3 >>
rect 3841 2513 3951 2567
<< via2 >>
rect 3848 2520 3944 2560
<< via1 >>
rect 3848 2520 3944 2560
<< m1 >>
rect 3265 513 3375 567
<< m2 >>
rect 3265 513 3375 567
<< via1 >>
rect 3272 520 3368 560
<< m1 >>
rect 3265 1713 3375 1767
<< m2 >>
rect 3265 1713 3375 1767
<< m3 >>
rect 3265 1713 3375 1767
<< via2 >>
rect 3272 1720 3368 1760
<< via1 >>
rect 3272 1720 3368 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< m3 >>
rect 3841 1713 3951 1767
<< via2 >>
rect 3848 1720 3944 1760
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< m3 >>
rect 3841 1713 3951 1767
<< via2 >>
rect 3848 1720 3944 1760
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< m3 >>
rect 3841 1713 3951 1767
<< via2 >>
rect 3848 1720 3944 1760
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< m3 >>
rect 3841 2113 3951 2167
<< via2 >>
rect 3848 2120 3944 2160
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< m3 >>
rect 3841 2113 3951 2167
<< via2 >>
rect 3848 2120 3944 2160
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< m3 >>
rect 3265 2113 3375 2167
<< via2 >>
rect 3272 2120 3368 2160
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< m3 >>
rect 3265 2113 3375 2167
<< via2 >>
rect 3272 2120 3368 2160
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< m3 >>
rect 3585 673 3631 727
<< via2 >>
rect 3592 680 3624 720
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< m3 >>
rect 3585 673 3631 727
<< via2 >>
rect 3592 680 3624 720
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< m3 >>
rect 3841 513 3951 567
<< via2 >>
rect 3848 520 3944 560
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< m3 >>
rect 3841 513 3951 567
<< via2 >>
rect 3848 520 3944 560
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3009 673 3055 727
<< m2 >>
rect 3009 673 3055 727
<< via1 >>
rect 3016 680 3048 720
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< m3 >>
rect 3073 1993 3183 2047
<< via2 >>
rect 3080 2000 3176 2040
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< m3 >>
rect 3649 1993 3759 2047
<< via2 >>
rect 3656 2000 3752 2040
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< m3 >>
rect 3649 2393 3759 2447
<< via2 >>
rect 3656 2400 3752 2440
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3073 2393 3183 2447
<< m2 >>
rect 3073 2393 3183 2447
<< via1 >>
rect 3080 2400 3176 2440
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< m3 >>
rect 3649 3193 3759 3247
<< via2 >>
rect 3656 3200 3752 3240
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3073 3193 3183 3247
<< m2 >>
rect 3073 3193 3183 3247
<< m3 >>
rect 3073 3193 3183 3247
<< via2 >>
rect 3080 3200 3176 3240
<< via1 >>
rect 3080 3200 3176 3240
<< m1 >>
rect 3073 3193 3183 3247
<< m2 >>
rect 3073 3193 3183 3247
<< via1 >>
rect 3080 3200 3176 3240
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< m3 >>
rect 3073 2793 3183 2847
<< via2 >>
rect 3080 2800 3176 2840
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< m3 >>
rect 3073 2793 3183 2847
<< via2 >>
rect 3080 2800 3176 2840
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< m3 >>
rect 3649 2793 3759 2847
<< via2 >>
rect 3656 2800 3752 2840
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3265 3313 3375 3367
<< m2 >>
rect 3265 3313 3375 3367
<< via1 >>
rect 3272 3320 3368 3360
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< m3 >>
rect 3009 3473 3055 3527
<< via2 >>
rect 3016 3480 3048 3520
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3585 3473 3631 3527
<< m2 >>
rect 3585 3473 3631 3527
<< via1 >>
rect 3592 3480 3624 3520
<< locali >>
rect 2203 1953 2361 2087
<< m1 >>
rect 2203 1953 2361 2087
<< m2 >>
rect 2203 1953 2361 2087
<< m3 >>
rect 2203 1953 2361 2087
<< via2 >>
rect 2210 1960 2354 2080
<< via1 >>
rect 2210 1960 2354 2080
<< viali >>
rect 2210 1960 2354 2080
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< m2 >>
rect 475 1953 633 2087
<< via1 >>
rect 482 1960 626 2080
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< m2 >>
rect 2203 3773 2361 3907
<< via1 >>
rect 2210 3780 2354 3900
<< viali >>
rect 2210 3780 2354 3900
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< m2 >>
rect 475 3773 633 3907
<< m3 >>
rect 475 3773 633 3907
<< via2 >>
rect 482 3780 626 3900
<< via1 >>
rect 482 3780 626 3900
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< m2 >>
rect 2203 5623 2361 5757
<< m3 >>
rect 2203 5623 2361 5757
<< via2 >>
rect 2210 5630 2354 5750
<< via1 >>
rect 2210 5630 2354 5750
<< viali >>
rect 2210 5630 2354 5750
<< m2 >>
rect 3463 1882 3606 1912
<< m3 >>
rect 3463 1882 3493 2312
<< m2 >>
rect 3463 2282 3621 2312
<< m3 >>
rect 3591 2282 3621 2312
<< m2 >>
rect 3015 2282 3621 2312
<< m3 >>
rect 3015 2282 3045 2312
<< m2 >>
rect 2887 2282 3045 2312
<< m3 >>
rect 2887 1882 2917 2312
<< m2 >>
rect 2887 1882 3030 1912
<< m1 >>
rect 3009 1873 3055 1927
<< m2 >>
rect 3009 1873 3055 1927
<< via1 >>
rect 3016 1880 3048 1920
<< m1 >>
rect 3585 1873 3631 1927
<< m2 >>
rect 3585 1873 3631 1927
<< via1 >>
rect 3592 1880 3624 1920
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3585 2273 3631 2327
<< m2 >>
rect 3585 2273 3631 2327
<< via1 >>
rect 3592 2280 3624 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< via1 >>
rect 3016 2280 3048 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< via1 >>
rect 3016 2280 3048 2320
<< m1 >>
rect 3009 2273 3055 2327
<< m2 >>
rect 3009 2273 3055 2327
<< via1 >>
rect 3016 2280 3048 2320
<< m2 >>
rect 3456 1875 3500 1919
<< m3 >>
rect 3456 1875 3500 1919
<< via2 >>
rect 3463 1882 3493 1912
<< m2 >>
rect 3456 2275 3500 2319
<< m3 >>
rect 3456 2275 3500 2319
<< via2 >>
rect 3463 2282 3493 2312
<< m2 >>
rect 3584 2275 3628 2319
<< m3 >>
rect 3584 2275 3628 2319
<< via2 >>
rect 3591 2282 3621 2312
<< m2 >>
rect 3584 2275 3628 2319
<< m3 >>
rect 3584 2275 3628 2319
<< via2 >>
rect 3591 2282 3621 2312
<< m2 >>
rect 3008 2275 3052 2319
<< m3 >>
rect 3008 2275 3052 2319
<< via2 >>
rect 3015 2282 3045 2312
<< m2 >>
rect 3008 2275 3052 2319
<< m3 >>
rect 3008 2275 3052 2319
<< via2 >>
rect 3015 2282 3045 2312
<< m2 >>
rect 2880 2275 2924 2319
<< m3 >>
rect 2880 2275 2924 2319
<< via2 >>
rect 2887 2282 2917 2312
<< m2 >>
rect 2880 1875 2924 1919
<< m3 >>
rect 2880 1875 2924 1919
<< via2 >>
rect 2887 1882 2917 1912
<< m2 >>
rect 2887 3082 3030 3112
<< m3 >>
rect 2887 2682 2917 3112
<< m2 >>
rect 2887 2682 3045 2712
<< m3 >>
rect 3015 2682 3045 2712
<< m2 >>
rect 3015 2682 3621 2712
<< m3 >>
rect 3591 2682 3621 2712
<< m2 >>
rect 3463 2682 3621 2712
<< m3 >>
rect 3463 2682 3493 3112
<< m2 >>
rect 3463 3082 3606 3112
<< m1 >>
rect 3585 3073 3631 3127
<< m2 >>
rect 3585 3073 3631 3127
<< via1 >>
rect 3592 3080 3624 3120
<< m1 >>
rect 3009 3073 3055 3127
<< m2 >>
rect 3009 3073 3055 3127
<< via1 >>
rect 3016 3080 3048 3120
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3009 2673 3055 2727
<< m2 >>
rect 3009 2673 3055 2727
<< via1 >>
rect 3016 2680 3048 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< via1 >>
rect 3592 2680 3624 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< via1 >>
rect 3592 2680 3624 2720
<< m1 >>
rect 3585 2673 3631 2727
<< m2 >>
rect 3585 2673 3631 2727
<< via1 >>
rect 3592 2680 3624 2720
<< m2 >>
rect 2880 3075 2924 3119
<< m3 >>
rect 2880 3075 2924 3119
<< via2 >>
rect 2887 3082 2917 3112
<< m2 >>
rect 2880 2675 2924 2719
<< m3 >>
rect 2880 2675 2924 2719
<< via2 >>
rect 2887 2682 2917 2712
<< m2 >>
rect 3008 2675 3052 2719
<< m3 >>
rect 3008 2675 3052 2719
<< via2 >>
rect 3015 2682 3045 2712
<< m2 >>
rect 3008 2675 3052 2719
<< m3 >>
rect 3008 2675 3052 2719
<< via2 >>
rect 3015 2682 3045 2712
<< m2 >>
rect 3584 2675 3628 2719
<< m3 >>
rect 3584 2675 3628 2719
<< via2 >>
rect 3591 2682 3621 2712
<< m2 >>
rect 3584 2675 3628 2719
<< m3 >>
rect 3584 2675 3628 2719
<< via2 >>
rect 3591 2682 3621 2712
<< m2 >>
rect 3456 2675 3500 2719
<< m3 >>
rect 3456 2675 3500 2719
<< via2 >>
rect 3463 2682 3493 2712
<< m2 >>
rect 3456 3075 3500 3119
<< m3 >>
rect 3456 3075 3500 3119
<< via2 >>
rect 3463 3082 3493 3112
<< m2 >>
rect 2791 523 3318 553
<< m3 >>
rect 2791 523 2821 2553
<< m2 >>
rect 2791 2523 3333 2553
<< m3 >>
rect 3303 2523 3333 2553
<< m3 >>
rect 3303 2523 3333 2953
<< m3 >>
rect 3303 2923 3333 2953
<< m2 >>
rect 3303 2923 3909 2953
<< m3 >>
rect 3879 2923 3909 2953
<< m3 >>
rect 3879 2538 3909 2953
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3841 2913 3951 2967
<< m2 >>
rect 3841 2913 3951 2967
<< via1 >>
rect 3848 2920 3944 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2913 3375 2967
<< m2 >>
rect 3265 2913 3375 2967
<< via1 >>
rect 3272 2920 3368 2960
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3265 2513 3375 2567
<< m2 >>
rect 3265 2513 3375 2567
<< via1 >>
rect 3272 2520 3368 2560
<< m1 >>
rect 3841 2513 3951 2567
<< m2 >>
rect 3841 2513 3951 2567
<< via1 >>
rect 3848 2520 3944 2560
<< m1 >>
rect 3265 513 3375 567
<< m2 >>
rect 3265 513 3375 567
<< via1 >>
rect 3272 520 3368 560
<< m2 >>
rect 2784 516 2828 560
<< m3 >>
rect 2784 516 2828 560
<< via2 >>
rect 2791 523 2821 553
<< m2 >>
rect 2784 2516 2828 2560
<< m3 >>
rect 2784 2516 2828 2560
<< via2 >>
rect 2791 2523 2821 2553
<< m2 >>
rect 3296 2516 3340 2560
<< m3 >>
rect 3296 2516 3340 2560
<< via2 >>
rect 3303 2523 3333 2553
<< m2 >>
rect 3296 2916 3340 2960
<< m3 >>
rect 3296 2916 3340 2960
<< via2 >>
rect 3303 2923 3333 2953
<< m2 >>
rect 3872 2916 3916 2960
<< m3 >>
rect 3872 2916 3916 2960
<< via2 >>
rect 3879 2923 3909 2953
<< m2 >>
rect 3031 683 3622 713
<< m3 >>
rect 3592 683 3622 713
<< m3 >>
rect 3592 523 3622 713
<< m2 >>
rect 3592 523 3910 553
<< m3 >>
rect 3880 523 3910 553
<< m3 >>
rect 3880 523 3910 1753
<< m3 >>
rect 3880 1723 3910 1753
<< m3 >>
rect 3880 1723 3910 2153
<< m3 >>
rect 3880 2123 3910 2153
<< m2 >>
rect 3304 2123 3910 2153
<< m3 >>
rect 3304 2123 3334 2153
<< m3 >>
rect 3304 1738 3334 2153
<< m1 >>
rect 3265 1713 3375 1767
<< m2 >>
rect 3265 1713 3375 1767
<< via1 >>
rect 3272 1720 3368 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 1713 3951 1767
<< m2 >>
rect 3841 1713 3951 1767
<< via1 >>
rect 3848 1720 3944 1760
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3841 2113 3951 2167
<< m2 >>
rect 3841 2113 3951 2167
<< via1 >>
rect 3848 2120 3944 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3265 2113 3375 2167
<< m2 >>
rect 3265 2113 3375 2167
<< via1 >>
rect 3272 2120 3368 2160
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3585 673 3631 727
<< m2 >>
rect 3585 673 3631 727
<< via1 >>
rect 3592 680 3624 720
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3841 513 3951 567
<< m2 >>
rect 3841 513 3951 567
<< via1 >>
rect 3848 520 3944 560
<< m1 >>
rect 3009 673 3055 727
<< m2 >>
rect 3009 673 3055 727
<< via1 >>
rect 3016 680 3048 720
<< m2 >>
rect 3585 676 3629 720
<< m3 >>
rect 3585 676 3629 720
<< via2 >>
rect 3592 683 3622 713
<< m2 >>
rect 3585 516 3629 560
<< m3 >>
rect 3585 516 3629 560
<< via2 >>
rect 3592 523 3622 553
<< m2 >>
rect 3873 516 3917 560
<< m3 >>
rect 3873 516 3917 560
<< via2 >>
rect 3880 523 3910 553
<< m2 >>
rect 3873 2116 3917 2160
<< m3 >>
rect 3873 2116 3917 2160
<< via2 >>
rect 3880 2123 3910 2153
<< m2 >>
rect 3297 2116 3341 2160
<< m3 >>
rect 3297 2116 3341 2160
<< via2 >>
rect 3304 2123 3334 2153
<< m2 >>
rect 3128 3317 3319 3347
<< m3 >>
rect 3128 2837 3158 3347
<< m2 >>
rect 3112 2837 3158 2867
<< m3 >>
rect 3112 2805 3142 2867
<< m2 >>
rect 3144 3205 3718 3235
<< m3 >>
rect 3688 3205 3718 3235
<< m2 >>
rect 3688 3205 4054 3235
<< m3 >>
rect 4024 2805 4054 3235
<< m2 >>
rect 3688 2805 4054 2835
<< m3 >>
rect 3688 2805 3718 2835
<< m2 >>
rect 3688 2805 4054 2835
<< m3 >>
rect 4024 2405 4054 2835
<< m2 >>
rect 3688 2405 4054 2435
<< m3 >>
rect 3688 2405 3718 2435
<< m2 >>
rect 3688 2405 4054 2435
<< m3 >>
rect 4024 2005 4054 2435
<< m2 >>
rect 3688 2005 4054 2035
<< m3 >>
rect 3688 2005 3718 2035
<< m2 >>
rect 3112 2005 3718 2035
<< m3 >>
rect 3112 2005 3142 2035
<< m2 >>
rect 2696 2005 3142 2035
<< m3 >>
rect 2696 2005 2726 2435
<< m2 >>
rect 2696 2405 3127 2435
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3073 1993 3183 2047
<< m2 >>
rect 3073 1993 3183 2047
<< via1 >>
rect 3080 2000 3176 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 1993 3759 2047
<< m2 >>
rect 3649 1993 3759 2047
<< via1 >>
rect 3656 2000 3752 2040
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3649 2393 3759 2447
<< m2 >>
rect 3649 2393 3759 2447
<< via1 >>
rect 3656 2400 3752 2440
<< m1 >>
rect 3073 2393 3183 2447
<< m2 >>
rect 3073 2393 3183 2447
<< via1 >>
rect 3080 2400 3176 2440
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3649 3193 3759 3247
<< m2 >>
rect 3649 3193 3759 3247
<< via1 >>
rect 3656 3200 3752 3240
<< m1 >>
rect 3073 3193 3183 3247
<< m2 >>
rect 3073 3193 3183 3247
<< via1 >>
rect 3080 3200 3176 3240
<< m1 >>
rect 3073 3193 3183 3247
<< m2 >>
rect 3073 3193 3183 3247
<< via1 >>
rect 3080 3200 3176 3240
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3073 2793 3183 2847
<< m2 >>
rect 3073 2793 3183 2847
<< via1 >>
rect 3080 2800 3176 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3649 2793 3759 2847
<< m2 >>
rect 3649 2793 3759 2847
<< via1 >>
rect 3656 2800 3752 2840
<< m1 >>
rect 3265 3313 3375 3367
<< m2 >>
rect 3265 3313 3375 3367
<< via1 >>
rect 3272 3320 3368 3360
<< m2 >>
rect 3121 3310 3165 3354
<< m3 >>
rect 3121 3310 3165 3354
<< via2 >>
rect 3128 3317 3158 3347
<< m2 >>
rect 3121 2830 3165 2874
<< m3 >>
rect 3121 2830 3165 2874
<< via2 >>
rect 3128 2837 3158 2867
<< m2 >>
rect 3105 2830 3149 2874
<< m3 >>
rect 3105 2830 3149 2874
<< via2 >>
rect 3112 2837 3142 2867
<< m2 >>
rect 3681 3198 3725 3242
<< m3 >>
rect 3681 3198 3725 3242
<< via2 >>
rect 3688 3205 3718 3235
<< m2 >>
rect 3681 3198 3725 3242
<< m3 >>
rect 3681 3198 3725 3242
<< via2 >>
rect 3688 3205 3718 3235
<< m2 >>
rect 4017 3198 4061 3242
<< m3 >>
rect 4017 3198 4061 3242
<< via2 >>
rect 4024 3205 4054 3235
<< m2 >>
rect 4017 2798 4061 2842
<< m3 >>
rect 4017 2798 4061 2842
<< via2 >>
rect 4024 2805 4054 2835
<< m2 >>
rect 3681 2798 3725 2842
<< m3 >>
rect 3681 2798 3725 2842
<< via2 >>
rect 3688 2805 3718 2835
<< m2 >>
rect 3681 2798 3725 2842
<< m3 >>
rect 3681 2798 3725 2842
<< via2 >>
rect 3688 2805 3718 2835
<< m2 >>
rect 4017 2798 4061 2842
<< m3 >>
rect 4017 2798 4061 2842
<< via2 >>
rect 4024 2805 4054 2835
<< m2 >>
rect 4017 2398 4061 2442
<< m3 >>
rect 4017 2398 4061 2442
<< via2 >>
rect 4024 2405 4054 2435
<< m2 >>
rect 3681 2398 3725 2442
<< m3 >>
rect 3681 2398 3725 2442
<< via2 >>
rect 3688 2405 3718 2435
<< m2 >>
rect 3681 2398 3725 2442
<< m3 >>
rect 3681 2398 3725 2442
<< via2 >>
rect 3688 2405 3718 2435
<< m2 >>
rect 4017 2398 4061 2442
<< m3 >>
rect 4017 2398 4061 2442
<< via2 >>
rect 4024 2405 4054 2435
<< m2 >>
rect 4017 1998 4061 2042
<< m3 >>
rect 4017 1998 4061 2042
<< via2 >>
rect 4024 2005 4054 2035
<< m2 >>
rect 3681 1998 3725 2042
<< m3 >>
rect 3681 1998 3725 2042
<< via2 >>
rect 3688 2005 3718 2035
<< m2 >>
rect 3681 1998 3725 2042
<< m3 >>
rect 3681 1998 3725 2042
<< via2 >>
rect 3688 2005 3718 2035
<< m2 >>
rect 3105 1998 3149 2042
<< m3 >>
rect 3105 1998 3149 2042
<< via2 >>
rect 3112 2005 3142 2035
<< m2 >>
rect 3105 1998 3149 2042
<< m3 >>
rect 3105 1998 3149 2042
<< via2 >>
rect 3112 2005 3142 2035
<< m2 >>
rect 2689 1998 2733 2042
<< m3 >>
rect 2689 1998 2733 2042
<< via2 >>
rect 2696 2005 2726 2035
<< m2 >>
rect 2689 2398 2733 2442
<< m3 >>
rect 2689 2398 2733 2442
<< via2 >>
rect 2696 2405 2726 2435
<< m3 >>
rect 2262 2024 2292 3511
<< m2 >>
rect 2262 3481 3044 3511
<< m3 >>
rect 3014 3481 3044 3511
<< m2 >>
rect 3014 3481 3605 3511
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3009 3473 3055 3527
<< m2 >>
rect 3009 3473 3055 3527
<< via1 >>
rect 3016 3480 3048 3520
<< m1 >>
rect 3585 3473 3631 3527
<< m2 >>
rect 3585 3473 3631 3527
<< via1 >>
rect 3592 3480 3624 3520
<< locali >>
rect 2203 1953 2361 2087
<< m1 >>
rect 2203 1953 2361 2087
<< viali >>
rect 2210 1960 2354 2080
<< m2 >>
rect 2255 3474 2299 3518
<< m3 >>
rect 2255 3474 2299 3518
<< via2 >>
rect 2262 3481 2292 3511
<< m2 >>
rect 3007 3474 3051 3518
<< m3 >>
rect 3007 3474 3051 3518
<< via2 >>
rect 3014 3481 3044 3511
<< m2 >>
rect 3007 3474 3051 3518
<< m3 >>
rect 3007 3474 3051 3518
<< via2 >>
rect 3014 3481 3044 3511
<< m2 >>
rect 549 2003 2100 2033
<< m3 >>
rect 2070 2003 2100 3857
<< m2 >>
rect 2070 3827 2277 3857
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< viali >>
rect 2210 3780 2354 3900
<< m2 >>
rect 2063 1996 2107 2040
<< m3 >>
rect 2063 1996 2107 2040
<< via2 >>
rect 2070 2003 2100 2033
<< m2 >>
rect 2063 3820 2107 3864
<< m3 >>
rect 2063 3820 2107 3864
<< via2 >>
rect 2070 3827 2100 3857
<< m3 >>
rect 534 3840 564 5503
<< m2 >>
rect 534 5473 2292 5503
<< m3 >>
rect 2262 5473 2292 5680
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< viali >>
rect 2210 5630 2354 5750
<< m2 >>
rect 527 5466 571 5510
<< m3 >>
rect 527 5466 571 5510
<< via2 >>
rect 534 5473 564 5503
<< m2 >>
rect 2255 5466 2299 5510
<< m3 >>
rect 2255 5466 2299 5510
<< via2 >>
rect 2262 5473 2292 5503
<< locali >>
rect 100 6240 4288 6290
<< locali >>
rect 100 100 4288 150
<< m1 >>
rect 100 150 150 6240
<< m1 >>
rect 4238 150 4288 6240
<< locali >>
rect 93 6233 157 6297
<< m1 >>
rect 93 6233 157 6297
<< viali >>
rect 100 6240 150 6290
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 4231 6233 4295 6297
<< m1 >>
rect 4231 6233 4295 6297
<< viali >>
rect 4238 6240 4288 6290
<< locali >>
rect 4231 93 4295 157
<< m1 >>
rect 4231 93 4295 157
<< viali >>
rect 4238 100 4288 150
<< locali >>
rect 0 6340 4388 6390
<< locali >>
rect 0 0 4388 50
<< m1 >>
rect 0 50 50 6340
<< m1 >>
rect 4338 50 4388 6340
<< locali >>
rect -7 6333 57 6397
<< m1 >>
rect -7 6333 57 6397
<< viali >>
rect 0 6340 50 6390
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 4331 6333 4395 6397
<< m1 >>
rect 4331 6333 4395 6397
<< viali >>
rect 4338 6340 4388 6390
<< locali >>
rect 4331 -7 4395 57
<< m1 >>
rect 4331 -7 4395 57
<< viali >>
rect 4338 0 4388 50
<< locali >>
rect 2888 3600 3176 3640
<< locali >>
rect 3464 3600 3752 3640
<< locali >>
rect 3848 3480 4008 3520
<< locali >>
rect 3464 800 3752 840
<< locali >>
rect 3848 680 4008 720
<< locali >>
rect 2888 800 3176 840
<< locali >>
rect 2936 1532 4288 1628
<< locali >>
rect 4231 1525 4295 1635
<< m1 >>
rect 4231 1525 4295 1635
<< viali >>
rect 4238 1532 4288 1628
<< locali >>
rect 2936 3772 4288 3868
<< locali >>
rect 4231 3765 4295 3875
<< m1 >>
rect 4231 3765 4295 3875
<< viali >>
rect 4238 3772 4288 3868
<< locali >>
rect 2936 972 4388 1068
<< locali >>
rect 4331 965 4395 1075
<< m1 >>
rect 4331 965 4395 1075
<< viali >>
rect 4338 972 4388 1068
<< locali >>
rect 2936 332 4388 428
<< locali >>
rect 4331 325 4395 435
<< m1 >>
rect 4331 325 4395 435
<< viali >>
rect 4338 332 4388 428
<< locali >>
rect 308 5630 626 5750
<< locali >>
rect 0 2164 2536 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 0 500 2536 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 0 3984 2536 4040
<< locali >>
rect -7 3977 57 4047
<< m1 >>
rect -7 3977 57 4047
<< viali >>
rect 0 3984 50 4040
<< locali >>
rect 0 2320 2536 2376
<< locali >>
rect -7 2313 57 2383
<< m1 >>
rect -7 2313 57 2383
<< viali >>
rect 0 2320 50 2376
<< locali >>
rect 0 5834 2536 5890
<< locali >>
rect -7 5827 57 5897
<< m1 >>
rect -7 5827 57 5897
<< viali >>
rect 0 5834 50 5890
<< locali >>
rect 0 4170 2536 4226
<< locali >>
rect -7 4163 57 4233
<< m1 >>
rect -7 4163 57 4233
<< viali >>
rect 0 4170 50 4226
<< labels >>
flabel m2 s 3463 1882 3606 1912 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 2887 3082 3030 3112 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 100 6240 4288 6290 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 0 6340 4388 6390 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m2 s 2791 523 3318 553 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
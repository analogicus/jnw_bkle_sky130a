magic
tech sky130A
magscale 1 2
timestamp 1744160456
<< metal4 >>
rect 0 0 1160 1160
rect 0 -225 1160 -200
rect 0 -475 126 -225
rect 1034 -475 1160 -225
rect 0 -525 1160 -475
<< via4 >>
rect 126 -475 1034 -225
<< mimcap2 >>
rect 80 1040 1080 1080
rect 80 120 120 1040
rect 1040 120 1080 1040
rect 80 80 1080 120
<< mimcap2contact >>
rect 120 120 1040 1040
<< metal5 >>
rect 96 1040 1064 1064
rect 96 120 120 1040
rect 1040 120 1064 1040
rect 96 -225 1064 120
rect 96 -475 126 -225
rect 1034 -475 1064 -225
rect 96 -500 1064 -475
<< labels >>
flabel metal4 s 0 0 1160 1160 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel metal4 s 0 -525 1160 -200 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 -525 1160 1160
<< end >>

magic
tech sky130A
magscale 1 1
timestamp 1748124392
<< checkpaint >>
rect 0 0 1 1
use JNWATR_NCH_4C5F0  diff1_MN1 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 904
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  diff1_MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 1304
box 0 0 576 240
use JNWATR_NCH_4C5F0  diff1_MN2 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 904
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  diff1_MN2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 1304
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP5 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 2804
box 0 0 576 240
use JNWATR_PCH_4CTAPBOT  load1_MP5_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 2164
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP6 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP6_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 2804
box 0 0 576 240
use JNWATR_PCH_4CTAPBOT  load1_MP6_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 2164
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP1 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  load1_MP1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 1764
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP2 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  load1_MP2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 1764
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN4 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN4_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN3 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN3_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN5 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 904
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 1304
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror1_MN5_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 292 0 1 664
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN6 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 904
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN6_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 1304
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror1_MN6_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 2020 0 1 664
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP3 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP3_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 868 0 1 2804
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP4 ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP4_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748124392
transform 1 0 1444 0 1 2804
box 0 0 576 240
<< m3 >>
rect 2387 936 2417 2440
<< m2 >>
rect 962 683 1538 713
<< m2 >>
rect 1396 2188 1539 2218
<< m3 >>
rect 1396 2188 1426 2618
<< m2 >>
rect 1396 2588 1554 2618
<< m2 >>
rect 1236 2588 1554 2618
<< m3 >>
rect 1236 2428 1266 2618
<< m3 >>
rect 1236 2188 1266 2458
<< m2 >>
rect 948 2188 1266 2218
<< m3 >>
rect 948 1420 978 2218
<< m2 >>
rect 948 1420 1266 1450
<< m3 >>
rect 1236 939 1266 1450
<< m2 >>
rect 1389 2181 1433 2225
<< m3 >>
rect 1389 2181 1433 2225
<< via2 >>
rect 1396 2188 1426 2218
<< m2 >>
rect 1389 2581 1433 2625
<< m3 >>
rect 1389 2581 1433 2625
<< via2 >>
rect 1396 2588 1426 2618
<< m2 >>
rect 1229 2581 1273 2625
<< m3 >>
rect 1229 2581 1273 2625
<< via2 >>
rect 1236 2588 1266 2618
<< m2 >>
rect 1229 2181 1273 2225
<< m3 >>
rect 1229 2181 1273 2225
<< via2 >>
rect 1236 2188 1266 2218
<< m2 >>
rect 941 2181 985 2225
<< m3 >>
rect 941 2181 985 2225
<< via2 >>
rect 948 2188 978 2218
<< m2 >>
rect 941 1413 985 1457
<< m3 >>
rect 941 1413 985 1457
<< via2 >>
rect 948 1420 978 1450
<< m2 >>
rect 1229 1413 1273 1457
<< m3 >>
rect 1229 1413 1273 1457
<< via2 >>
rect 1236 1420 1266 1450
<< m2 >>
rect 1827 520 1986 550
<< m3 >>
rect 1956 520 1986 1238
<< m2 >>
rect 1620 1208 1986 1238
<< m2 >>
rect 1059 1208 1650 1238
<< m2 >>
rect 1949 513 1993 557
<< m3 >>
rect 1949 513 1993 557
<< via2 >>
rect 1956 520 1986 550
<< m2 >>
rect 1949 1201 1993 1245
<< m3 >>
rect 1949 1201 1993 1245
<< via2 >>
rect 1956 1208 1986 1238
<< m2 >>
rect 387 2588 978 2618
<< m2 >>
rect 820 2588 978 2618
<< m3 >>
rect 820 2588 850 2826
<< m2 >>
rect 820 2796 2002 2826
<< m3 >>
rect 1972 2588 2002 2826
<< m2 >>
rect 1972 2588 2130 2618
<< m2 >>
rect 1812 2588 2130 2618
<< m3 >>
rect 1812 2428 1842 2618
<< m2 >>
rect 1812 2428 1986 2458
<< m3 >>
rect 1956 1372 1986 2458
<< m2 >>
rect 1812 1372 1986 1402
<< m3 >>
rect 1812 939 1842 1402
<< m2 >>
rect 813 2581 857 2625
<< m3 >>
rect 813 2581 857 2625
<< via2 >>
rect 820 2588 850 2618
<< m2 >>
rect 813 2789 857 2833
<< m3 >>
rect 813 2789 857 2833
<< via2 >>
rect 820 2796 850 2826
<< m2 >>
rect 1965 2789 2009 2833
<< m3 >>
rect 1965 2789 2009 2833
<< via2 >>
rect 1972 2796 2002 2826
<< m2 >>
rect 1965 2581 2009 2625
<< m3 >>
rect 1965 2581 2009 2625
<< via2 >>
rect 1972 2588 2002 2618
<< m2 >>
rect 1805 2581 1849 2625
<< m3 >>
rect 1805 2581 1849 2625
<< via2 >>
rect 1812 2588 1842 2618
<< m2 >>
rect 1805 2421 1849 2465
<< m3 >>
rect 1805 2421 1849 2465
<< via2 >>
rect 1812 2428 1842 2458
<< m2 >>
rect 1949 2421 1993 2465
<< m3 >>
rect 1949 2421 1993 2465
<< via2 >>
rect 1956 2428 1986 2458
<< m2 >>
rect 1949 1365 1993 1409
<< m3 >>
rect 1949 1365 1993 1409
<< via2 >>
rect 1956 1372 1986 1402
<< m2 >>
rect 1805 1365 1849 1409
<< m3 >>
rect 1805 1365 1849 1409
<< via2 >>
rect 1812 1372 1842 1402
<< m3 >>
rect 2100 1068 2130 1099
<< m2 >>
rect 1636 1068 2130 1098
<< m3 >>
rect 1636 940 1666 1098
<< m2 >>
rect 1380 940 1666 970
<< m3 >>
rect 1380 940 1410 1098
<< m2 >>
rect 1076 1068 1410 1098
<< m3 >>
rect 1076 940 1106 1098
<< m2 >>
rect 836 940 1106 970
<< m3 >>
rect 836 940 866 1114
<< m2 >>
rect 372 1084 866 1114
<< m2 >>
rect 372 1084 754 1114
<< m3 >>
rect 724 1084 754 2058
<< m2 >>
rect 724 2028 1251 2058
<< m2 >>
rect 2093 1061 2137 1105
<< m3 >>
rect 2093 1061 2137 1105
<< via2 >>
rect 2100 1068 2130 1098
<< m2 >>
rect 1629 1061 1673 1105
<< m3 >>
rect 1629 1061 1673 1105
<< via2 >>
rect 1636 1068 1666 1098
<< m2 >>
rect 1629 933 1673 977
<< m3 >>
rect 1629 933 1673 977
<< via2 >>
rect 1636 940 1666 970
<< m2 >>
rect 1373 933 1417 977
<< m3 >>
rect 1373 933 1417 977
<< via2 >>
rect 1380 940 1410 970
<< m2 >>
rect 1373 1061 1417 1105
<< m3 >>
rect 1373 1061 1417 1105
<< via2 >>
rect 1380 1068 1410 1098
<< m2 >>
rect 1069 1061 1113 1105
<< m3 >>
rect 1069 1061 1113 1105
<< via2 >>
rect 1076 1068 1106 1098
<< m2 >>
rect 1069 933 1113 977
<< m3 >>
rect 1069 933 1113 977
<< via2 >>
rect 1076 940 1106 970
<< m2 >>
rect 829 933 873 977
<< m3 >>
rect 829 933 873 977
<< via2 >>
rect 836 940 866 970
<< m2 >>
rect 829 1077 873 1121
<< m3 >>
rect 829 1077 873 1121
<< via2 >>
rect 836 1084 866 1114
<< m2 >>
rect 717 1077 761 1121
<< m3 >>
rect 717 1077 761 1121
<< via2 >>
rect 724 1084 754 1114
<< m2 >>
rect 717 2021 761 2065
<< m3 >>
rect 717 2021 761 2065
<< via2 >>
rect 724 2028 754 2058
<< locali >>
rect 100 3158 2788 3208
<< locali >>
rect 100 100 2788 150
<< m1 >>
rect 100 150 150 3158
<< m1 >>
rect 2738 150 2788 3158
<< locali >>
rect 93 3151 157 3215
<< m1 >>
rect 93 3151 157 3215
<< viali >>
rect 100 3158 150 3208
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2731 3151 2795 3215
<< m1 >>
rect 2731 3151 2795 3215
<< viali >>
rect 2738 3158 2788 3208
<< locali >>
rect 2731 93 2795 157
<< m1 >>
rect 2731 93 2795 157
<< viali >>
rect 2738 100 2788 150
<< locali >>
rect 0 3258 2888 3308
<< locali >>
rect 0 0 2888 50
<< m1 >>
rect 0 50 50 3258
<< m1 >>
rect 2838 50 2888 3258
<< locali >>
rect -7 3251 57 3315
<< m1 >>
rect -7 3251 57 3315
<< viali >>
rect 0 3258 50 3308
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2831 3251 2895 3315
<< m1 >>
rect 2831 3251 2895 3315
<< viali >>
rect 2838 3258 2888 3308
<< locali >>
rect 2831 -7 2895 57
<< m1 >>
rect 2831 -7 2895 57
<< viali >>
rect 2838 0 2888 50
<< locali >>
rect 244 2704 532 2744
<< locali >>
rect 628 2584 788 2624
<< locali >>
rect 1972 2704 2260 2744
<< locali >>
rect 820 2304 1108 2344
<< locali >>
rect 1396 2304 1684 2344
<< locali >>
rect 1780 2184 1940 2224
<< locali >>
rect 1396 804 1684 844
<< locali >>
rect 820 804 1108 844
<< locali >>
rect 1204 684 1364 724
<< locali >>
rect 244 1204 532 1244
<< locali >>
rect 628 1084 788 1124
<< locali >>
rect 1972 1204 2260 1244
<< locali >>
rect 820 2704 1108 2744
<< locali >>
rect 1396 2704 1684 2744
<< locali >>
rect 100 1376 2788 1472
<< locali >>
rect 93 1369 157 1479
<< m1 >>
rect 93 1369 157 1479
<< viali >>
rect 100 1376 150 1472
<< locali >>
rect 2731 1369 2795 1479
<< m1 >>
rect 2731 1369 2795 1479
<< viali >>
rect 2738 1376 2788 1472
<< locali >>
rect 0 2876 2888 2972
<< locali >>
rect -7 2869 57 2979
<< m1 >>
rect -7 2869 57 2979
<< viali >>
rect 0 2876 50 2972
<< locali >>
rect 2831 2869 2895 2979
<< m1 >>
rect 2831 2869 2895 2979
<< viali >>
rect 2838 2876 2888 2972
<< locali >>
rect 0 1836 2888 1932
<< locali >>
rect -7 1829 57 1939
<< m1 >>
rect -7 1829 57 1939
<< viali >>
rect 0 1836 50 1932
<< locali >>
rect 2831 1829 2895 1939
<< m1 >>
rect 2831 1829 2895 1939
<< viali >>
rect 2838 1836 2888 1932
<< locali >>
rect 100 336 2788 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< locali >>
rect 2731 329 2795 439
<< m1 >>
rect 2731 329 2795 439
<< viali >>
rect 2738 336 2788 432
<< m1 >>
rect 2349 2417 2459 2471
<< m2 >>
rect 2349 2417 2459 2471
<< m3 >>
rect 2349 2417 2459 2471
<< via2 >>
rect 2356 2424 2452 2464
<< via1 >>
rect 2356 2424 2452 2464
<< m1 >>
rect 2349 917 2459 971
<< m2 >>
rect 2349 917 2459 971
<< m3 >>
rect 2349 917 2459 971
<< via2 >>
rect 2356 924 2452 964
<< via1 >>
rect 2356 924 2452 964
<< m1 >>
rect 1517 677 1563 731
<< m2 >>
rect 1517 677 1563 731
<< via1 >>
rect 1524 684 1556 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 1197 917 1307 971
<< m2 >>
rect 1197 917 1307 971
<< m3 >>
rect 1197 917 1307 971
<< via2 >>
rect 1204 924 1300 964
<< via1 >>
rect 1204 924 1300 964
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< m3 >>
rect 941 2177 987 2231
<< via2 >>
rect 948 2184 980 2224
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 1517 2177 1563 2231
<< m2 >>
rect 1517 2177 1563 2231
<< via1 >>
rect 1524 2184 1556 2224
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< m3 >>
rect 1197 2417 1307 2471
<< via2 >>
rect 1204 2424 1300 2464
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< m3 >>
rect 1197 2417 1307 2471
<< via2 >>
rect 1204 2424 1300 2464
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1517 2577 1563 2631
<< m2 >>
rect 1517 2577 1563 2631
<< via1 >>
rect 1524 2584 1556 2624
<< m1 >>
rect 1517 2577 1563 2631
<< m2 >>
rect 1517 2577 1563 2631
<< via1 >>
rect 1524 2584 1556 2624
<< m1 >>
rect 1005 1197 1115 1251
<< m2 >>
rect 1005 1197 1115 1251
<< via1 >>
rect 1012 1204 1108 1244
<< m1 >>
rect 1581 1197 1691 1251
<< m2 >>
rect 1581 1197 1691 1251
<< via1 >>
rect 1588 1204 1684 1244
<< m1 >>
rect 1581 1197 1691 1251
<< m2 >>
rect 1581 1197 1691 1251
<< via1 >>
rect 1588 1204 1684 1244
<< m1 >>
rect 1773 517 1883 571
<< m2 >>
rect 1773 517 1883 571
<< via1 >>
rect 1780 524 1876 564
<< m1 >>
rect 1773 917 1883 971
<< m2 >>
rect 1773 917 1883 971
<< m3 >>
rect 1773 917 1883 971
<< via2 >>
rect 1780 924 1876 964
<< via1 >>
rect 1780 924 1876 964
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 2093 2577 2139 2631
<< m2 >>
rect 2093 2577 2139 2631
<< via1 >>
rect 2100 2584 2132 2624
<< m1 >>
rect 2093 2577 2139 2631
<< m2 >>
rect 2093 2577 2139 2631
<< via1 >>
rect 2100 2584 2132 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 1773 2417 1883 2471
<< m2 >>
rect 1773 2417 1883 2471
<< m3 >>
rect 1773 2417 1883 2471
<< via2 >>
rect 1780 2424 1876 2464
<< via1 >>
rect 1780 2424 1876 2464
<< m1 >>
rect 1773 2417 1883 2471
<< m2 >>
rect 1773 2417 1883 2471
<< via1 >>
rect 1780 2424 1876 2464
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 365 1077 411 1131
<< m2 >>
rect 365 1077 411 1131
<< via1 >>
rect 372 1084 404 1124
<< m1 >>
rect 365 1077 411 1131
<< m2 >>
rect 365 1077 411 1131
<< via1 >>
rect 372 1084 404 1124
<< m1 >>
rect 2093 1077 2139 1131
<< m2 >>
rect 2093 1077 2139 1131
<< m3 >>
rect 2093 1077 2139 1131
<< via2 >>
rect 2100 1084 2132 1124
<< via1 >>
rect 2100 1084 2132 1124
<< m1 >>
rect 2093 1077 2139 1131
<< m2 >>
rect 2093 1077 2139 1131
<< via1 >>
rect 2100 1084 2132 1124
<< labels >>
flabel locali s 100 3158 2788 3208 0 FreeSans 400 0 0 0 VSS
port 4 nsew signal bidirectional
flabel locali s 0 3258 2888 3308 0 FreeSans 400 0 0 0 VDD
port 5 nsew signal bidirectional
flabel m1 s 948 1084 980 1124 0 FreeSans 400 0 0 0 VIP
port 6 nsew signal bidirectional
flabel m1 s 1524 1084 1556 1124 0 FreeSans 400 0 0 0 VIN
port 7 nsew signal bidirectional
flabel m3 s 2387 936 2417 2440 0 FreeSans 400 0 0 0 VO
port 8 nsew signal bidirectional
flabel m2 s 962 683 1538 713 0 FreeSans 400 0 0 0 I_BIAS
port 9 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1746404937
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 1464
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 1464
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 2904
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 2904
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 2504
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 2504
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 3304
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 3704
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 3304
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 3704
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 264
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1610 0 1 200
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1610 0 1 3740
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1610 0 1 1970
box 0 0 2236 1720
<< m1 >>
rect 849 1877 895 1931
<< m2 >>
rect 849 1877 895 1931
<< via1 >>
rect 856 1884 888 1924
<< m1 >>
rect 273 1877 319 1931
<< m2 >>
rect 273 1877 319 1931
<< via1 >>
rect 280 1884 312 1924
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< m3 >>
rect 273 2277 319 2331
<< via2 >>
rect 280 2284 312 2324
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< via1 >>
rect 856 2284 888 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< m3 >>
rect 849 2277 895 2331
<< via2 >>
rect 856 2284 888 2324
<< via1 >>
rect 856 2284 888 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< via1 >>
rect 856 2284 888 2324
<< m1 >>
rect 849 3077 895 3131
<< m2 >>
rect 849 3077 895 3131
<< via1 >>
rect 856 3084 888 3124
<< m1 >>
rect 273 3077 319 3131
<< m2 >>
rect 273 3077 319 3131
<< via1 >>
rect 280 3084 312 3124
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< m3 >>
rect 849 2677 895 2731
<< via2 >>
rect 856 2684 888 2724
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< via1 >>
rect 280 2684 312 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< m3 >>
rect 273 2677 319 2731
<< via2 >>
rect 280 2684 312 2724
<< via1 >>
rect 280 2684 312 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< via1 >>
rect 280 2684 312 2724
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< m3 >>
rect 1105 2917 1215 2971
<< via2 >>
rect 1112 2924 1208 2964
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< m3 >>
rect 1105 2917 1215 2971
<< via2 >>
rect 1112 2924 1208 2964
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< m3 >>
rect 529 2917 639 2971
<< via2 >>
rect 536 2924 632 2964
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< m3 >>
rect 529 2917 639 2971
<< via2 >>
rect 536 2924 632 2964
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 1105 2517 1215 2571
<< m2 >>
rect 1105 2517 1215 2571
<< m3 >>
rect 1105 2517 1215 2571
<< via2 >>
rect 1112 2524 1208 2564
<< via1 >>
rect 1112 2524 1208 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< m3 >>
rect 529 2517 639 2571
<< via2 >>
rect 536 2524 632 2564
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< m3 >>
rect 529 2517 639 2571
<< via2 >>
rect 536 2524 632 2564
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 517 639 571
<< m2 >>
rect 529 517 639 571
<< via1 >>
rect 536 524 632 564
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< m3 >>
rect 1105 1717 1215 1771
<< via2 >>
rect 1112 1724 1208 1764
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< m3 >>
rect 1105 1717 1215 1771
<< via2 >>
rect 1112 1724 1208 1764
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< m3 >>
rect 1105 1717 1215 1771
<< via2 >>
rect 1112 1724 1208 1764
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 529 1717 639 1771
<< m2 >>
rect 529 1717 639 1771
<< m3 >>
rect 529 1717 639 1771
<< via2 >>
rect 536 1724 632 1764
<< via1 >>
rect 536 1724 632 1764
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< m3 >>
rect 529 2117 639 2171
<< via2 >>
rect 536 2124 632 2164
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< m3 >>
rect 529 2117 639 2171
<< via2 >>
rect 536 2124 632 2164
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< m3 >>
rect 1105 2117 1215 2171
<< via2 >>
rect 1112 2124 1208 2164
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< m3 >>
rect 1105 2117 1215 2171
<< via2 >>
rect 1112 2124 1208 2164
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< m3 >>
rect 849 677 895 731
<< via2 >>
rect 856 684 888 724
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< m3 >>
rect 849 677 895 731
<< via2 >>
rect 856 684 888 724
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< m3 >>
rect 1105 517 1215 571
<< via2 >>
rect 1112 524 1208 564
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< m3 >>
rect 1105 517 1215 571
<< via2 >>
rect 1112 524 1208 564
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 273 677 319 731
<< m2 >>
rect 273 677 319 731
<< via1 >>
rect 280 684 312 724
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< m3 >>
rect 913 1997 1023 2051
<< via2 >>
rect 920 2004 1016 2044
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< m3 >>
rect 337 1997 447 2051
<< via2 >>
rect 344 2004 440 2044
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< m3 >>
rect 337 2397 447 2451
<< via2 >>
rect 344 2404 440 2444
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 913 2397 1023 2451
<< m2 >>
rect 913 2397 1023 2451
<< via1 >>
rect 920 2404 1016 2444
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< m3 >>
rect 913 3197 1023 3251
<< via2 >>
rect 920 3204 1016 3244
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< m3 >>
rect 337 3197 447 3251
<< via2 >>
rect 344 3204 440 3244
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 913 2797 1023 2851
<< m2 >>
rect 913 2797 1023 2851
<< via1 >>
rect 920 2804 1016 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< m3 >>
rect 337 2797 447 2851
<< via2 >>
rect 344 2804 440 2844
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 1105 3317 1215 3371
<< m2 >>
rect 1105 3317 1215 3371
<< via1 >>
rect 1112 3324 1208 3364
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< m3 >>
rect 849 3477 895 3531
<< via2 >>
rect 856 3484 888 3524
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< m3 >>
rect 849 3477 895 3531
<< via2 >>
rect 856 3484 888 3524
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 529 3317 639 3371
<< m2 >>
rect 529 3317 639 3371
<< via1 >>
rect 536 3324 632 3364
<< locali >>
rect 3513 1653 3671 1787
<< m1 >>
rect 3513 1653 3671 1787
<< m2 >>
rect 3513 1653 3671 1787
<< m3 >>
rect 3513 1653 3671 1787
<< via2 >>
rect 3520 1660 3664 1780
<< via1 >>
rect 3520 1660 3664 1780
<< viali >>
rect 3520 1660 3664 1780
<< locali >>
rect 1785 1653 1943 1787
<< m1 >>
rect 1785 1653 1943 1787
<< m2 >>
rect 1785 1653 1943 1787
<< via1 >>
rect 1792 1660 1936 1780
<< viali >>
rect 1792 1660 1936 1780
<< locali >>
rect 3513 5193 3671 5327
<< m1 >>
rect 3513 5193 3671 5327
<< m2 >>
rect 3513 5193 3671 5327
<< via1 >>
rect 3520 5200 3664 5320
<< viali >>
rect 3520 5200 3664 5320
<< locali >>
rect 1785 5193 1943 5327
<< m1 >>
rect 1785 5193 1943 5327
<< m2 >>
rect 1785 5193 1943 5327
<< via1 >>
rect 1792 5200 1936 5320
<< viali >>
rect 1792 5200 1936 5320
<< locali >>
rect 3513 3423 3671 3557
<< m1 >>
rect 3513 3423 3671 3557
<< m2 >>
rect 3513 3423 3671 3557
<< via1 >>
rect 3520 3430 3664 3550
<< viali >>
rect 3520 3430 3664 3550
<< m2 >>
rect 150 1886 293 1916
<< m3 >>
rect 150 1886 180 2316
<< m2 >>
rect 150 2286 308 2316
<< m3 >>
rect 278 2286 308 2316
<< m2 >>
rect 278 2286 884 2316
<< m3 >>
rect 854 2286 884 2316
<< m2 >>
rect 726 2286 884 2316
<< m3 >>
rect 726 1886 756 2316
<< m2 >>
rect 726 1886 869 1916
<< m1 >>
rect 849 1877 895 1931
<< m2 >>
rect 849 1877 895 1931
<< via1 >>
rect 856 1884 888 1924
<< m1 >>
rect 273 1877 319 1931
<< m2 >>
rect 273 1877 319 1931
<< via1 >>
rect 280 1884 312 1924
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 273 2277 319 2331
<< m2 >>
rect 273 2277 319 2331
<< via1 >>
rect 280 2284 312 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< via1 >>
rect 856 2284 888 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< via1 >>
rect 856 2284 888 2324
<< m1 >>
rect 849 2277 895 2331
<< m2 >>
rect 849 2277 895 2331
<< via1 >>
rect 856 2284 888 2324
<< m2 >>
rect 143 1879 187 1923
<< m3 >>
rect 143 1879 187 1923
<< via2 >>
rect 150 1886 180 1916
<< m2 >>
rect 143 2279 187 2323
<< m3 >>
rect 143 2279 187 2323
<< via2 >>
rect 150 2286 180 2316
<< m2 >>
rect 271 2279 315 2323
<< m3 >>
rect 271 2279 315 2323
<< via2 >>
rect 278 2286 308 2316
<< m2 >>
rect 271 2279 315 2323
<< m3 >>
rect 271 2279 315 2323
<< via2 >>
rect 278 2286 308 2316
<< m2 >>
rect 847 2279 891 2323
<< m3 >>
rect 847 2279 891 2323
<< via2 >>
rect 854 2286 884 2316
<< m2 >>
rect 847 2279 891 2323
<< m3 >>
rect 847 2279 891 2323
<< via2 >>
rect 854 2286 884 2316
<< m2 >>
rect 719 2279 763 2323
<< m3 >>
rect 719 2279 763 2323
<< via2 >>
rect 726 2286 756 2316
<< m2 >>
rect 719 1879 763 1923
<< m3 >>
rect 719 1879 763 1923
<< via2 >>
rect 726 1886 756 1916
<< m2 >>
rect 150 3086 293 3116
<< m3 >>
rect 150 2686 180 3116
<< m2 >>
rect 150 2686 308 2716
<< m3 >>
rect 278 2686 308 2716
<< m2 >>
rect 278 2686 884 2716
<< m3 >>
rect 854 2686 884 2716
<< m2 >>
rect 726 2686 884 2716
<< m3 >>
rect 726 2686 756 3116
<< m2 >>
rect 726 3086 869 3116
<< m1 >>
rect 849 3077 895 3131
<< m2 >>
rect 849 3077 895 3131
<< via1 >>
rect 856 3084 888 3124
<< m1 >>
rect 273 3077 319 3131
<< m2 >>
rect 273 3077 319 3131
<< via1 >>
rect 280 3084 312 3124
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 849 2677 895 2731
<< m2 >>
rect 849 2677 895 2731
<< via1 >>
rect 856 2684 888 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< via1 >>
rect 280 2684 312 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< via1 >>
rect 280 2684 312 2724
<< m1 >>
rect 273 2677 319 2731
<< m2 >>
rect 273 2677 319 2731
<< via1 >>
rect 280 2684 312 2724
<< m2 >>
rect 143 3079 187 3123
<< m3 >>
rect 143 3079 187 3123
<< via2 >>
rect 150 3086 180 3116
<< m2 >>
rect 143 2679 187 2723
<< m3 >>
rect 143 2679 187 2723
<< via2 >>
rect 150 2686 180 2716
<< m2 >>
rect 271 2679 315 2723
<< m3 >>
rect 271 2679 315 2723
<< via2 >>
rect 278 2686 308 2716
<< m2 >>
rect 271 2679 315 2723
<< m3 >>
rect 271 2679 315 2723
<< via2 >>
rect 278 2686 308 2716
<< m2 >>
rect 847 2679 891 2723
<< m3 >>
rect 847 2679 891 2723
<< via2 >>
rect 854 2686 884 2716
<< m2 >>
rect 847 2679 891 2723
<< m3 >>
rect 847 2679 891 2723
<< via2 >>
rect 854 2686 884 2716
<< m2 >>
rect 719 2679 763 2723
<< m3 >>
rect 719 2679 763 2723
<< via2 >>
rect 726 2686 756 2716
<< m2 >>
rect 719 3079 763 3123
<< m3 >>
rect 719 3079 763 3123
<< via2 >>
rect 726 3086 756 3116
<< m2 >>
rect 55 527 582 557
<< m3 >>
rect 55 527 85 2557
<< m2 >>
rect 55 2527 597 2557
<< m3 >>
rect 567 2527 597 2557
<< m3 >>
rect 567 2527 597 2957
<< m3 >>
rect 567 2927 597 2957
<< m2 >>
rect 567 2927 1173 2957
<< m3 >>
rect 1143 2927 1173 2957
<< m3 >>
rect 1143 2542 1173 2957
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 1105 2917 1215 2971
<< m2 >>
rect 1105 2917 1215 2971
<< via1 >>
rect 1112 2924 1208 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 529 2917 639 2971
<< m2 >>
rect 529 2917 639 2971
<< via1 >>
rect 536 2924 632 2964
<< m1 >>
rect 1105 2517 1215 2571
<< m2 >>
rect 1105 2517 1215 2571
<< via1 >>
rect 1112 2524 1208 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 2517 639 2571
<< m2 >>
rect 529 2517 639 2571
<< via1 >>
rect 536 2524 632 2564
<< m1 >>
rect 529 517 639 571
<< m2 >>
rect 529 517 639 571
<< via1 >>
rect 536 524 632 564
<< m2 >>
rect 48 520 92 564
<< m3 >>
rect 48 520 92 564
<< via2 >>
rect 55 527 85 557
<< m2 >>
rect 48 2520 92 2564
<< m3 >>
rect 48 2520 92 2564
<< via2 >>
rect 55 2527 85 2557
<< m2 >>
rect 560 2520 604 2564
<< m3 >>
rect 560 2520 604 2564
<< via2 >>
rect 567 2527 597 2557
<< m2 >>
rect 560 2920 604 2964
<< m3 >>
rect 560 2920 604 2964
<< via2 >>
rect 567 2927 597 2957
<< m2 >>
rect 1136 2920 1180 2964
<< m3 >>
rect 1136 2920 1180 2964
<< via2 >>
rect 1143 2927 1173 2957
<< m2 >>
rect 294 687 885 717
<< m3 >>
rect 855 687 885 717
<< m3 >>
rect 855 527 885 717
<< m2 >>
rect 855 527 1173 557
<< m3 >>
rect 1143 527 1173 557
<< m3 >>
rect 1143 527 1173 1757
<< m3 >>
rect 1143 1727 1173 1757
<< m3 >>
rect 1143 1727 1173 2157
<< m3 >>
rect 1143 2127 1173 2157
<< m2 >>
rect 567 2127 1173 2157
<< m3 >>
rect 567 2127 597 2157
<< m3 >>
rect 567 1742 597 2157
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 1105 1717 1215 1771
<< m2 >>
rect 1105 1717 1215 1771
<< via1 >>
rect 1112 1724 1208 1764
<< m1 >>
rect 529 1717 639 1771
<< m2 >>
rect 529 1717 639 1771
<< via1 >>
rect 536 1724 632 1764
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 529 2117 639 2171
<< m2 >>
rect 529 2117 639 2171
<< via1 >>
rect 536 2124 632 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 1105 2117 1215 2171
<< m2 >>
rect 1105 2117 1215 2171
<< via1 >>
rect 1112 2124 1208 2164
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 849 677 895 731
<< m2 >>
rect 849 677 895 731
<< via1 >>
rect 856 684 888 724
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 1105 517 1215 571
<< m2 >>
rect 1105 517 1215 571
<< via1 >>
rect 1112 524 1208 564
<< m1 >>
rect 273 677 319 731
<< m2 >>
rect 273 677 319 731
<< via1 >>
rect 280 684 312 724
<< m2 >>
rect 848 680 892 724
<< m3 >>
rect 848 680 892 724
<< via2 >>
rect 855 687 885 717
<< m2 >>
rect 848 520 892 564
<< m3 >>
rect 848 520 892 564
<< via2 >>
rect 855 527 885 557
<< m2 >>
rect 1136 520 1180 564
<< m3 >>
rect 1136 520 1180 564
<< via2 >>
rect 1143 527 1173 557
<< m2 >>
rect 1136 2120 1180 2164
<< m3 >>
rect 1136 2120 1180 2164
<< via2 >>
rect 1143 2127 1173 2157
<< m2 >>
rect 560 2120 604 2164
<< m3 >>
rect 560 2120 604 2164
<< via2 >>
rect 567 2127 597 2157
<< m2 >>
rect 1159 3321 1318 3351
<< m3 >>
rect 1288 2809 1318 3351
<< m2 >>
rect 952 2809 1318 2839
<< m2 >>
rect 952 3209 1302 3239
<< m3 >>
rect 952 3209 982 3239
<< m2 >>
rect 376 3209 982 3239
<< m3 >>
rect 376 3209 406 3239
<< m2 >>
rect 56 3209 406 3239
<< m3 >>
rect 56 2809 86 3239
<< m2 >>
rect 56 2809 406 2839
<< m3 >>
rect 376 2809 406 2839
<< m2 >>
rect -40 2809 406 2839
<< m3 >>
rect -40 2409 -10 2839
<< m2 >>
rect -40 2409 406 2439
<< m3 >>
rect 376 2409 406 2439
<< m2 >>
rect -40 2409 406 2439
<< m3 >>
rect -40 2009 -10 2439
<< m2 >>
rect -40 2009 406 2039
<< m3 >>
rect 376 2009 406 2039
<< m2 >>
rect 376 2009 982 2039
<< m3 >>
rect 952 2009 982 2039
<< m2 >>
rect 952 2009 1318 2039
<< m3 >>
rect 1288 2009 1318 2439
<< m2 >>
rect 967 2409 1318 2439
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 913 1997 1023 2051
<< m2 >>
rect 913 1997 1023 2051
<< via1 >>
rect 920 2004 1016 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 1997 447 2051
<< m2 >>
rect 337 1997 447 2051
<< via1 >>
rect 344 2004 440 2044
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 337 2397 447 2451
<< m2 >>
rect 337 2397 447 2451
<< via1 >>
rect 344 2404 440 2444
<< m1 >>
rect 913 2397 1023 2451
<< m2 >>
rect 913 2397 1023 2451
<< via1 >>
rect 920 2404 1016 2444
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 913 3197 1023 3251
<< m2 >>
rect 913 3197 1023 3251
<< via1 >>
rect 920 3204 1016 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 337 3197 447 3251
<< m2 >>
rect 337 3197 447 3251
<< via1 >>
rect 344 3204 440 3244
<< m1 >>
rect 913 2797 1023 2851
<< m2 >>
rect 913 2797 1023 2851
<< via1 >>
rect 920 2804 1016 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 337 2797 447 2851
<< m2 >>
rect 337 2797 447 2851
<< via1 >>
rect 344 2804 440 2844
<< m1 >>
rect 1105 3317 1215 3371
<< m2 >>
rect 1105 3317 1215 3371
<< via1 >>
rect 1112 3324 1208 3364
<< m2 >>
rect 1281 3314 1325 3358
<< m3 >>
rect 1281 3314 1325 3358
<< via2 >>
rect 1288 3321 1318 3351
<< m2 >>
rect 1281 2802 1325 2846
<< m3 >>
rect 1281 2802 1325 2846
<< via2 >>
rect 1288 2809 1318 2839
<< m2 >>
rect 945 3202 989 3246
<< m3 >>
rect 945 3202 989 3246
<< via2 >>
rect 952 3209 982 3239
<< m2 >>
rect 945 3202 989 3246
<< m3 >>
rect 945 3202 989 3246
<< via2 >>
rect 952 3209 982 3239
<< m2 >>
rect 369 3202 413 3246
<< m3 >>
rect 369 3202 413 3246
<< via2 >>
rect 376 3209 406 3239
<< m2 >>
rect 369 3202 413 3246
<< m3 >>
rect 369 3202 413 3246
<< via2 >>
rect 376 3209 406 3239
<< m2 >>
rect 49 3202 93 3246
<< m3 >>
rect 49 3202 93 3246
<< via2 >>
rect 56 3209 86 3239
<< m2 >>
rect 49 2802 93 2846
<< m3 >>
rect 49 2802 93 2846
<< via2 >>
rect 56 2809 86 2839
<< m2 >>
rect 369 2802 413 2846
<< m3 >>
rect 369 2802 413 2846
<< via2 >>
rect 376 2809 406 2839
<< m2 >>
rect 369 2802 413 2846
<< m3 >>
rect 369 2802 413 2846
<< via2 >>
rect 376 2809 406 2839
<< m2 >>
rect -47 2802 -3 2846
<< m3 >>
rect -47 2802 -3 2846
<< via2 >>
rect -40 2809 -10 2839
<< m2 >>
rect -47 2402 -3 2446
<< m3 >>
rect -47 2402 -3 2446
<< via2 >>
rect -40 2409 -10 2439
<< m2 >>
rect 369 2402 413 2446
<< m3 >>
rect 369 2402 413 2446
<< via2 >>
rect 376 2409 406 2439
<< m2 >>
rect 369 2402 413 2446
<< m3 >>
rect 369 2402 413 2446
<< via2 >>
rect 376 2409 406 2439
<< m2 >>
rect -47 2402 -3 2446
<< m3 >>
rect -47 2402 -3 2446
<< via2 >>
rect -40 2409 -10 2439
<< m2 >>
rect -47 2002 -3 2046
<< m3 >>
rect -47 2002 -3 2046
<< via2 >>
rect -40 2009 -10 2039
<< m2 >>
rect 369 2002 413 2046
<< m3 >>
rect 369 2002 413 2046
<< via2 >>
rect 376 2009 406 2039
<< m2 >>
rect 369 2002 413 2046
<< m3 >>
rect 369 2002 413 2046
<< via2 >>
rect 376 2009 406 2039
<< m2 >>
rect 945 2002 989 2046
<< m3 >>
rect 945 2002 989 2046
<< via2 >>
rect 952 2009 982 2039
<< m2 >>
rect 945 2002 989 2046
<< m3 >>
rect 945 2002 989 2046
<< via2 >>
rect 952 2009 982 2039
<< m2 >>
rect 1281 2002 1325 2046
<< m3 >>
rect 1281 2002 1325 2046
<< via2 >>
rect 1288 2009 1318 2039
<< m2 >>
rect 1281 2402 1325 2446
<< m3 >>
rect 1281 2402 1325 2446
<< via2 >>
rect 1288 2409 1318 2439
<< m3 >>
rect 3573 1724 3603 3307
<< m2 >>
rect 1717 3277 3603 3307
<< m3 >>
rect 1717 3277 1747 3515
<< m2 >>
rect 853 3485 1747 3515
<< m3 >>
rect 853 3485 883 3515
<< m3 >>
rect 853 3325 883 3515
<< m2 >>
rect 580 3325 883 3355
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 849 3477 895 3531
<< m2 >>
rect 849 3477 895 3531
<< via1 >>
rect 856 3484 888 3524
<< m1 >>
rect 529 3317 639 3371
<< m2 >>
rect 529 3317 639 3371
<< via1 >>
rect 536 3324 632 3364
<< locali >>
rect 3513 1653 3671 1787
<< m1 >>
rect 3513 1653 3671 1787
<< viali >>
rect 3520 1660 3664 1780
<< m2 >>
rect 3566 3270 3610 3314
<< m3 >>
rect 3566 3270 3610 3314
<< via2 >>
rect 3573 3277 3603 3307
<< m2 >>
rect 1710 3270 1754 3314
<< m3 >>
rect 1710 3270 1754 3314
<< via2 >>
rect 1717 3277 1747 3307
<< m2 >>
rect 1710 3478 1754 3522
<< m3 >>
rect 1710 3478 1754 3522
<< via2 >>
rect 1717 3485 1747 3515
<< m2 >>
rect 846 3478 890 3522
<< m3 >>
rect 846 3478 890 3522
<< via2 >>
rect 853 3485 883 3515
<< m2 >>
rect 846 3318 890 3362
<< m3 >>
rect 846 3318 890 3362
<< via2 >>
rect 853 3325 883 3355
<< m2 >>
rect 1858 1703 3473 1733
<< m3 >>
rect 3443 1703 3473 5269
<< m2 >>
rect 3443 5239 3586 5269
<< locali >>
rect 1785 1653 1943 1787
<< m1 >>
rect 1785 1653 1943 1787
<< viali >>
rect 1792 1660 1936 1780
<< locali >>
rect 3513 5193 3671 5327
<< m1 >>
rect 3513 5193 3671 5327
<< viali >>
rect 3520 5200 3664 5320
<< m2 >>
rect 3436 1696 3480 1740
<< m3 >>
rect 3436 1696 3480 1740
<< via2 >>
rect 3443 1703 3473 1733
<< m2 >>
rect 3436 5232 3480 5276
<< m3 >>
rect 3436 5232 3480 5276
<< via2 >>
rect 3443 5239 3473 5269
<< m2 >>
rect 1858 5241 3169 5271
<< m3 >>
rect 3139 3465 3169 5271
<< m2 >>
rect 3139 3465 3586 3495
<< locali >>
rect 1785 5193 1943 5327
<< m1 >>
rect 1785 5193 1943 5327
<< viali >>
rect 1792 5200 1936 5320
<< locali >>
rect 3513 3423 3671 3557
<< m1 >>
rect 3513 3423 3671 3557
<< viali >>
rect 3520 3430 3664 3550
<< m2 >>
rect 3132 5234 3176 5278
<< m3 >>
rect 3132 5234 3176 5278
<< via2 >>
rect 3139 5241 3169 5271
<< m2 >>
rect 3132 3458 3176 3502
<< m3 >>
rect 3132 3458 3176 3502
<< via2 >>
rect 3139 3465 3169 3495
<< locali >>
rect 100 5510 3946 5560
<< locali >>
rect 100 100 3946 150
<< m1 >>
rect 100 150 150 5510
<< m1 >>
rect 3896 150 3946 5510
<< locali >>
rect 93 5503 157 5567
<< m1 >>
rect 93 5503 157 5567
<< viali >>
rect 100 5510 150 5560
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 3889 5503 3953 5567
<< m1 >>
rect 3889 5503 3953 5567
<< viali >>
rect 3896 5510 3946 5560
<< locali >>
rect 3889 93 3953 157
<< m1 >>
rect 3889 93 3953 157
<< viali >>
rect 3896 100 3946 150
<< locali >>
rect 0 5610 4046 5660
<< locali >>
rect 0 0 4046 50
<< m1 >>
rect 0 50 50 5610
<< m1 >>
rect 3996 50 4046 5610
<< locali >>
rect -7 5603 57 5667
<< m1 >>
rect -7 5603 57 5667
<< viali >>
rect 0 5610 50 5660
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 3989 5603 4053 5667
<< m1 >>
rect 3989 5603 4053 5667
<< viali >>
rect 3996 5610 4046 5660
<< locali >>
rect 3989 -7 4053 57
<< m1 >>
rect 3989 -7 4053 57
<< viali >>
rect 3996 0 4046 50
<< locali >>
rect 1618 3430 1936 3550
<< locali >>
rect 1610 1864 3946 1920
<< locali >>
rect 3889 1857 3953 1927
<< m1 >>
rect 3889 1857 3953 1927
<< viali >>
rect 3896 1864 3946 1920
<< locali >>
rect 1610 200 3946 256
<< locali >>
rect 3889 193 3953 263
<< m1 >>
rect 3889 193 3953 263
<< viali >>
rect 3896 200 3946 256
<< locali >>
rect 1610 5404 3946 5460
<< locali >>
rect 3889 5397 3953 5467
<< m1 >>
rect 3889 5397 3953 5467
<< viali >>
rect 3896 5404 3946 5460
<< locali >>
rect 1610 3740 3946 3796
<< locali >>
rect 3889 3733 3953 3803
<< m1 >>
rect 3889 3733 3953 3803
<< viali >>
rect 3896 3740 3946 3796
<< locali >>
rect 1610 3634 3946 3690
<< locali >>
rect 3889 3627 3953 3697
<< m1 >>
rect 3889 3627 3953 3697
<< viali >>
rect 3896 3634 3946 3690
<< locali >>
rect 1610 1970 3946 2026
<< locali >>
rect 3889 1963 3953 2033
<< m1 >>
rect 3889 1963 3953 2033
<< viali >>
rect 3896 1970 3946 2026
<< locali >>
rect 728 3604 1016 3644
<< locali >>
rect 152 3604 440 3644
<< locali >>
rect 536 3484 696 3524
<< locali >>
rect 728 804 1016 844
<< locali >>
rect 1112 684 1272 724
<< locali >>
rect 152 804 440 844
<< locali >>
rect 0 1536 1352 1632
<< locali >>
rect -7 1529 57 1639
<< m1 >>
rect -7 1529 57 1639
<< viali >>
rect 0 1536 50 1632
<< locali >>
rect 0 3776 1352 3872
<< locali >>
rect -7 3769 57 3879
<< m1 >>
rect -7 3769 57 3879
<< viali >>
rect 0 3776 50 3872
<< locali >>
rect 100 976 1352 1072
<< locali >>
rect 93 969 157 1079
<< m1 >>
rect 93 969 157 1079
<< viali >>
rect 100 976 150 1072
<< locali >>
rect 100 336 1352 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< labels >>
flabel m2 s 150 1886 293 1916 0 FreeSans 400 0 0 0 IN+
port 14 nsew signal bidirectional
flabel m2 s 150 3086 293 3116 0 FreeSans 400 0 0 0 IN-
port 15 nsew signal bidirectional
flabel locali s 0 5610 4046 5660 0 FreeSans 400 0 0 0 VDD
port 16 nsew signal bidirectional
flabel locali s 100 5510 3946 5560 0 FreeSans 400 0 0 0 VSS
port 17 nsew signal bidirectional
flabel m2 s 55 527 582 557 0 FreeSans 400 0 0 0 OUT
port 18 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1746190069
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 5710 5908 5760
<< locali >>
rect -100 -100 5908 -50
<< m1 >>
rect -100 -50 -50 5710
<< m1 >>
rect 5858 -50 5908 5710
<< locali >>
rect -107 5703 -43 5767
<< m1 >>
rect -107 5703 -43 5767
<< viali >>
rect -100 5710 -50 5760
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 5851 5703 5915 5767
<< m1 >>
rect 5851 5703 5915 5767
<< viali >>
rect 5858 5710 5908 5760
<< locali >>
rect 5851 -107 5915 -43
<< m1 >>
rect 5851 -107 5915 -43
<< viali >>
rect 5858 -100 5908 -50
<< locali >>
rect -200 5810 6008 5860
<< locali >>
rect -200 -200 6008 -150
<< m1 >>
rect -200 -150 -150 5810
<< m1 >>
rect 5958 -150 6008 5810
<< locali >>
rect -207 5803 -143 5867
<< m1 >>
rect -207 5803 -143 5867
<< viali >>
rect -200 5810 -150 5860
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 5951 5803 6015 5867
<< m1 >>
rect 5951 5803 6015 5867
<< viali >>
rect 5958 5810 6008 5860
<< locali >>
rect 5951 -207 6015 -143
<< m1 >>
rect 5951 -207 6015 -143
<< viali >>
rect 5958 -200 6008 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 5858 5710
<< labels >>
flabel locali s -100 5710 5908 5760 0 FreeSans 400 0 0 0 VDD
port 57 nsew signal bidirectional
flabel locali s -200 5810 6008 5860 0 FreeSans 400 0 0 0 VSS
port 58 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1748249007
<< checkpaint >>
rect 0 0 1 1
use JNWTR_RPPO4  res_RH2 ../JNW_TR_SKY130A
timestamp 1748249007
transform 1 0 200 0 1 3074
box 0 0 940 1720
use JNWTR_RPPO4  res_RH3 ../JNW_TR_SKY130A
timestamp 1748249007
transform 1 0 200 0 1 1304
box 0 0 940 1720
use JNWTR_RPPO4  res_RH1 ../JNW_TR_SKY130A
timestamp 1748249007
transform 1 0 200 0 1 4844
box 0 0 940 1720
use AALMISC_CAP50f  CM1 ../AAL_MISC_SKY130A
timestamp 1748249007
transform 1 0 200 0 1 6764
box 0 0 580 842
use JNWATR_NCH_2C1F2  MN1 ../JNW_ATR_SKY130A
timestamp 1748249007
transform 1 0 292 0 1 504
box 0 0 512 400
use JNWATR_NCH_2CTAPTOP  MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748249007
transform 1 0 292 0 1 904
box 0 0 512 240
use JNWATR_NCH_2CTAPBOT  MN1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748249007
transform 1 0 292 0 1 264
box 0 0 512 240
<< m2 >>
rect 453 4572 692 4602
<< m3 >>
rect 662 4572 692 6378
<< m2 >>
rect 662 6348 885 6378
<< m2 >>
rect 655 4565 699 4609
<< m3 >>
rect 655 4565 699 4609
<< via2 >>
rect 662 4572 692 4602
<< m2 >>
rect 655 6341 699 6385
<< m3 >>
rect 655 6341 699 6385
<< via2 >>
rect 662 6348 692 6378
<< m3 >>
rect 870 2972 900 4587
<< m2 >>
rect 438 2972 900 3002
<< m3 >>
rect 438 2827 468 3002
<< m2 >>
rect 863 2965 907 3009
<< m3 >>
rect 863 2965 907 3009
<< via2 >>
rect 870 2972 900 3002
<< m2 >>
rect 431 2965 475 3009
<< m3 >>
rect 431 2965 475 3009
<< via2 >>
rect 438 2972 468 3002
<< m2 >>
rect 264 6807 487 6837
<< m3 >>
rect 264 519 294 6837
<< m2 >>
rect 264 519 615 549
<< m2 >>
rect 257 6800 301 6844
<< m3 >>
rect 257 6800 301 6844
<< via2 >>
rect 264 6807 294 6837
<< m2 >>
rect 257 512 301 556
<< m3 >>
rect 257 512 301 556
<< via2 >>
rect 264 519 294 549
<< locali >>
rect 100 7656 1240 7706
<< locali >>
rect 100 100 1240 150
<< m1 >>
rect 100 150 150 7656
<< m1 >>
rect 1190 150 1240 7656
<< locali >>
rect 93 7649 157 7713
<< m1 >>
rect 93 7649 157 7713
<< viali >>
rect 100 7656 150 7706
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1183 7649 1247 7713
<< m1 >>
rect 1183 7649 1247 7713
<< viali >>
rect 1190 7656 1240 7706
<< locali >>
rect 1183 93 1247 157
<< m1 >>
rect 1183 93 1247 157
<< viali >>
rect 1190 100 1240 150
<< locali >>
rect 0 7756 1340 7806
<< locali >>
rect 0 0 1340 50
<< m1 >>
rect 0 50 50 7756
<< m1 >>
rect 1290 50 1340 7756
<< locali >>
rect -7 7749 57 7813
<< m1 >>
rect -7 7749 57 7813
<< viali >>
rect 0 7756 50 7806
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1283 7749 1347 7813
<< m1 >>
rect 1283 7749 1347 7813
<< viali >>
rect 1290 7756 1340 7806
<< locali >>
rect 1283 -7 1347 57
<< m1 >>
rect 1283 -7 1347 57
<< viali >>
rect 1290 0 1340 50
<< locali >>
rect 814 2764 1132 2884
<< locali >>
rect 100 4738 1240 4794
<< locali >>
rect 93 4731 157 4801
<< m1 >>
rect 93 4731 157 4801
<< viali >>
rect 100 4738 150 4794
<< locali >>
rect 1183 4731 1247 4801
<< m1 >>
rect 1183 4731 1247 4801
<< viali >>
rect 1190 4738 1240 4794
<< locali >>
rect 100 3074 1240 3130
<< locali >>
rect 93 3067 157 3137
<< m1 >>
rect 93 3067 157 3137
<< viali >>
rect 100 3074 150 3130
<< locali >>
rect 1183 3067 1247 3137
<< m1 >>
rect 1183 3067 1247 3137
<< viali >>
rect 1190 3074 1240 3130
<< locali >>
rect 100 2968 1240 3024
<< locali >>
rect 93 2961 157 3031
<< m1 >>
rect 93 2961 157 3031
<< viali >>
rect 100 2968 150 3024
<< locali >>
rect 1183 2961 1247 3031
<< m1 >>
rect 1183 2961 1247 3031
<< viali >>
rect 1190 2968 1240 3024
<< locali >>
rect 100 1304 1240 1360
<< locali >>
rect 93 1297 157 1367
<< m1 >>
rect 93 1297 157 1367
<< viali >>
rect 100 1304 150 1360
<< locali >>
rect 1183 1297 1247 1367
<< m1 >>
rect 1183 1297 1247 1367
<< viali >>
rect 1190 1304 1240 1360
<< locali >>
rect 100 6508 1240 6564
<< locali >>
rect 93 6501 157 6571
<< m1 >>
rect 93 6501 157 6571
<< viali >>
rect 100 6508 150 6564
<< locali >>
rect 1183 6501 1247 6571
<< m1 >>
rect 1183 6501 1247 6571
<< viali >>
rect 1190 6508 1240 6564
<< locali >>
rect 100 4844 1240 4900
<< locali >>
rect 93 4837 157 4907
<< m1 >>
rect 93 4837 157 4907
<< viali >>
rect 100 4844 150 4900
<< locali >>
rect 1183 4837 1247 4907
<< m1 >>
rect 1183 4837 1247 4907
<< viali >>
rect 1190 4844 1240 4900
<< locali >>
rect 244 804 532 844
<< locali >>
rect 100 976 1240 1072
<< locali >>
rect 93 969 157 1079
<< m1 >>
rect 93 969 157 1079
<< viali >>
rect 100 976 150 1072
<< locali >>
rect 1183 969 1247 1079
<< m1 >>
rect 1183 969 1247 1079
<< viali >>
rect 1190 976 1240 1072
<< locali >>
rect 100 336 1240 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< locali >>
rect 1183 329 1247 439
<< m1 >>
rect 1183 329 1247 439
<< viali >>
rect 1190 336 1240 432
<< locali >>
rect 100 7016 1240 7045
<< locali >>
rect 193 7009 787 7052
<< m1 >>
rect 193 7009 787 7052
<< m2 >>
rect 193 7009 787 7052
<< m3 >>
rect 193 7009 787 7052
<< viali >>
rect 200 7016 780 7045
<< via1 >>
rect 200 7016 780 7045
<< via2 >>
rect 200 7016 780 7045
<< locali >>
rect 93 7009 157 7052
<< m1 >>
rect 93 7009 157 7052
<< viali >>
rect 100 7016 150 7045
<< locali >>
rect 1183 7009 1247 7052
<< m1 >>
rect 1183 7009 1247 7052
<< viali >>
rect 1190 7016 1240 7045
<< locali >>
rect 375 4527 533 4661
<< m1 >>
rect 375 4527 533 4661
<< m2 >>
rect 375 4527 533 4661
<< via1 >>
rect 382 4534 526 4654
<< viali >>
rect 382 4534 526 4654
<< locali >>
rect 807 6297 965 6431
<< m1 >>
rect 807 6297 965 6431
<< m2 >>
rect 807 6297 965 6431
<< via1 >>
rect 814 6304 958 6424
<< viali >>
rect 814 6304 958 6424
<< locali >>
rect 807 4527 965 4661
<< m1 >>
rect 807 4527 965 4661
<< m2 >>
rect 807 4527 965 4661
<< m3 >>
rect 807 4527 965 4661
<< via2 >>
rect 814 4534 958 4654
<< via1 >>
rect 814 4534 958 4654
<< viali >>
rect 814 4534 958 4654
<< locali >>
rect 375 2757 533 2891
<< m1 >>
rect 375 2757 533 2891
<< m2 >>
rect 375 2757 533 2891
<< m3 >>
rect 375 2757 533 2891
<< via2 >>
rect 382 2764 526 2884
<< via1 >>
rect 382 2764 526 2884
<< viali >>
rect 382 2764 526 2884
<< m1 >>
rect 557 517 667 571
<< m2 >>
rect 557 517 667 571
<< via1 >>
rect 564 524 660 564
use single_stage_OTA U2_single_stage_OTA 
transform 1 0 1390 0 1 0
box 0 0 2686 9614
use temp_affected_current U1_temp_affected_current 
transform 1 0 4076 0 1 0
box 0 0 1890 10704
<< labels >>
flabel locali s 0 7756 1340 7806 0 FreeSans 400 0 0 0 VDD
port 4 nsew signal bidirectional
flabel locali s 100 7656 1240 7706 0 FreeSans 400 0 0 0 VSS
port 5 nsew signal bidirectional
flabel m1 s 372 684 404 724 0 FreeSans 400 0 0 0 reset
port 7 nsew signal bidirectional
<< properties >>
<< end >>

magic
tech sky130A
magscale 1 1
timestamp 1748204603
<< checkpaint >>
rect 0 0 1 1
use JNWATR_NCH_4C5F0  diff1_MN1 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 548 0 1 904
box 0 0 576 400
use JNWATR_NCH_4C5F0  diff1_MN2 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 904
box 0 0 576 400
use JNWATR_PCH_12C5F0  load1_MP5 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 2804
box 0 0 832 400
use JNWATR_PCH_12C5F0  load1_MP6 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2804
box 0 0 832 400
use JNWATR_PCH_12C5F0  load1_MP1 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 3204
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP  load1_MP1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 3604
box 0 0 832 240
use JNWATR_PCH_12C5F0  load1_MP2 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 3204
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP  load1_MP2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 3604
box 0 0 832 240
use JNWATR_NCH_4C5F0  mirror2_MN4 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN4_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN3 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 548 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN3_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 548 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN5 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 548 0 1 1304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 548 0 1 1704
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN6 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 1304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN6_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 1704
box 0 0 576 240
use JNWATR_PCH_12C5F0  load1_MP3 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2404
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT  load1_MP3_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2164
box 0 0 832 240
use JNWATR_PCH_12C5F0  load1_MP4 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 2404
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT  load1_MP4_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 1124 0 1 2164
box 0 0 832 240
<< m2 >>
rect 930 2825 1521 2855
<< m3 >>
rect 1491 1336 1521 2855
<< m2 >>
rect 1484 2818 1528 2862
<< m3 >>
rect 1484 2818 1528 2862
<< via2 >>
rect 1491 2825 1521 2855
<< m2 >>
rect 642 683 1218 713
<< m2 >>
rect 387 3388 1234 3418
<< m2 >>
rect 1076 3388 1234 3418
<< m3 >>
rect 1076 2588 1106 3418
<< m2 >>
rect 1076 2588 1234 2618
<< m2 >>
rect 916 2588 1234 2618
<< m3 >>
rect 916 2428 946 2618
<< m2 >>
rect 916 2428 1090 2458
<< m3 >>
rect 1060 924 1090 2458
<< m2 >>
rect 931 924 1090 954
<< m2 >>
rect 1069 3381 1113 3425
<< m3 >>
rect 1069 3381 1113 3425
<< via2 >>
rect 1076 3388 1106 3418
<< m2 >>
rect 1069 2581 1113 2625
<< m3 >>
rect 1069 2581 1113 2625
<< via2 >>
rect 1076 2588 1106 2618
<< m2 >>
rect 909 2581 953 2625
<< m3 >>
rect 909 2581 953 2625
<< via2 >>
rect 916 2588 946 2618
<< m2 >>
rect 909 2421 953 2465
<< m3 >>
rect 909 2421 953 2465
<< via2 >>
rect 916 2428 946 2458
<< m2 >>
rect 1053 2421 1097 2465
<< m3 >>
rect 1053 2421 1097 2465
<< via2 >>
rect 1060 2428 1090 2458
<< m2 >>
rect 1053 917 1097 961
<< m3 >>
rect 1053 917 1097 961
<< via2 >>
rect 1060 924 1090 954
<< m2 >>
rect 1507 520 1666 550
<< m3 >>
rect 1636 520 1666 1238
<< m2 >>
rect 1300 1208 1666 1238
<< m2 >>
rect 739 1208 1330 1238
<< m2 >>
rect 1629 513 1673 557
<< m3 >>
rect 1629 513 1673 557
<< via2 >>
rect 1636 520 1666 550
<< m2 >>
rect 1629 1201 1673 1245
<< m3 >>
rect 1629 1201 1673 1245
<< via2 >>
rect 1636 1208 1666 1238
<< m2 >>
rect 244 2588 387 2618
<< m3 >>
rect 244 2588 274 3018
<< m2 >>
rect 244 2988 402 3018
<< m2 >>
rect 372 2988 1234 3018
<< m2 >>
rect 1204 2988 1634 3018
<< m3 >>
rect 1604 2428 1634 3018
<< m2 >>
rect 1604 2428 1778 2458
<< m3 >>
rect 1748 924 1778 2458
<< m2 >>
rect 1507 924 1778 954
<< m2 >>
rect 237 2581 281 2625
<< m3 >>
rect 237 2581 281 2625
<< via2 >>
rect 244 2588 274 2618
<< m2 >>
rect 237 2981 281 3025
<< m3 >>
rect 237 2981 281 3025
<< via2 >>
rect 244 2988 274 3018
<< m2 >>
rect 1597 2981 1641 3025
<< m3 >>
rect 1597 2981 1641 3025
<< via2 >>
rect 1604 2988 1634 3018
<< m2 >>
rect 1597 2421 1641 2465
<< m3 >>
rect 1597 2421 1641 2465
<< via2 >>
rect 1604 2428 1634 2458
<< m2 >>
rect 1741 2421 1785 2465
<< m3 >>
rect 1741 2421 1785 2465
<< via2 >>
rect 1748 2428 1778 2458
<< m2 >>
rect 1741 917 1785 961
<< m3 >>
rect 1741 917 1785 961
<< via2 >>
rect 1748 924 1778 954
<< m2 >>
rect 628 1484 1219 1514
<< m2 >>
rect 500 1484 658 1514
<< m3 >>
rect 500 1484 530 2522
<< m2 >>
rect 500 2492 706 2522
<< m3 >>
rect 676 2492 706 3258
<< m2 >>
rect 676 3228 931 3258
<< m2 >>
rect 493 1477 537 1521
<< m3 >>
rect 493 1477 537 1521
<< via2 >>
rect 500 1484 530 1514
<< m2 >>
rect 493 2485 537 2529
<< m3 >>
rect 493 2485 537 2529
<< via2 >>
rect 500 2492 530 2522
<< m2 >>
rect 669 2485 713 2529
<< m3 >>
rect 669 2485 713 2529
<< via2 >>
rect 676 2492 706 2522
<< m2 >>
rect 669 3221 713 3265
<< m3 >>
rect 669 3221 713 3265
<< via2 >>
rect 676 3228 706 3258
<< locali >>
rect 100 3958 2148 4008
<< locali >>
rect 100 100 2148 150
<< m1 >>
rect 100 150 150 3958
<< m1 >>
rect 2098 150 2148 3958
<< locali >>
rect 93 3951 157 4015
<< m1 >>
rect 93 3951 157 4015
<< viali >>
rect 100 3958 150 4008
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2091 3951 2155 4015
<< m1 >>
rect 2091 3951 2155 4015
<< viali >>
rect 2098 3958 2148 4008
<< locali >>
rect 2091 93 2155 157
<< m1 >>
rect 2091 93 2155 157
<< viali >>
rect 2098 100 2148 150
<< locali >>
rect 0 4058 2248 4108
<< locali >>
rect 0 0 2248 50
<< m1 >>
rect 0 50 50 4058
<< m1 >>
rect 2198 50 2248 4058
<< locali >>
rect -7 4051 57 4115
<< m1 >>
rect -7 4051 57 4115
<< viali >>
rect 0 4058 50 4108
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2191 4051 2255 4115
<< m1 >>
rect 2191 4051 2255 4115
<< viali >>
rect 2198 4058 2248 4108
<< locali >>
rect 2191 -7 2255 57
<< m1 >>
rect 2191 -7 2255 57
<< viali >>
rect 2198 0 2248 50
<< locali >>
rect 1076 3104 1364 3144
<< locali >>
rect 1716 2984 1876 3024
<< locali >>
rect 244 3104 532 3144
<< locali >>
rect 244 3504 532 3544
<< locali >>
rect 1076 3504 1364 3544
<< locali >>
rect 1716 3384 1876 3424
<< locali >>
rect 1076 804 1364 844
<< locali >>
rect 500 804 788 844
<< locali >>
rect 884 684 1044 724
<< locali >>
rect 500 1604 788 1644
<< locali >>
rect 884 1484 1044 1524
<< locali >>
rect 1076 1604 1364 1644
<< locali >>
rect 244 2704 532 2744
<< locali >>
rect 1076 2704 1364 2744
<< locali >>
rect 0 3676 2248 3772
<< locali >>
rect -7 3669 57 3779
<< m1 >>
rect -7 3669 57 3779
<< viali >>
rect 0 3676 50 3772
<< locali >>
rect 2191 3669 2255 3779
<< m1 >>
rect 2191 3669 2255 3779
<< viali >>
rect 2198 3676 2248 3772
<< locali >>
rect 100 336 2148 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< locali >>
rect 2091 329 2155 439
<< m1 >>
rect 2091 329 2155 439
<< viali >>
rect 2098 336 2148 432
<< locali >>
rect 100 1776 2148 1872
<< locali >>
rect 93 1769 157 1879
<< m1 >>
rect 93 1769 157 1879
<< viali >>
rect 100 1776 150 1872
<< locali >>
rect 2091 1769 2155 1879
<< m1 >>
rect 2091 1769 2155 1879
<< viali >>
rect 2098 1776 2148 1872
<< locali >>
rect 0 2236 2248 2332
<< locali >>
rect -7 2229 57 2339
<< m1 >>
rect -7 2229 57 2339
<< viali >>
rect 0 2236 50 2332
<< locali >>
rect 2191 2229 2255 2339
<< m1 >>
rect 2191 2229 2255 2339
<< viali >>
rect 2198 2236 2248 2332
<< m1 >>
rect 877 2817 987 2871
<< m2 >>
rect 877 2817 987 2871
<< via1 >>
rect 884 2824 980 2864
<< m1 >>
rect 1453 1317 1563 1371
<< m2 >>
rect 1453 1317 1563 1371
<< m3 >>
rect 1453 1317 1563 1371
<< via2 >>
rect 1460 1324 1556 1364
<< via1 >>
rect 1460 1324 1556 1364
<< m1 >>
rect 1197 677 1243 731
<< m2 >>
rect 1197 677 1243 731
<< via1 >>
rect 1204 684 1236 724
<< m1 >>
rect 621 677 667 731
<< m2 >>
rect 621 677 667 731
<< via1 >>
rect 628 684 660 724
<< m1 >>
rect 877 917 987 971
<< m2 >>
rect 877 917 987 971
<< via1 >>
rect 884 924 980 964
<< m1 >>
rect 365 3377 411 3431
<< m2 >>
rect 365 3377 411 3431
<< via1 >>
rect 372 3384 404 3424
<< m1 >>
rect 1197 3377 1243 3431
<< m2 >>
rect 1197 3377 1243 3431
<< via1 >>
rect 1204 3384 1236 3424
<< m1 >>
rect 1197 3377 1243 3431
<< m2 >>
rect 1197 3377 1243 3431
<< via1 >>
rect 1204 3384 1236 3424
<< m1 >>
rect 877 2417 987 2471
<< m2 >>
rect 877 2417 987 2471
<< m3 >>
rect 877 2417 987 2471
<< via2 >>
rect 884 2424 980 2464
<< via1 >>
rect 884 2424 980 2464
<< m1 >>
rect 877 2417 987 2471
<< m2 >>
rect 877 2417 987 2471
<< via1 >>
rect 884 2424 980 2464
<< m1 >>
rect 1197 2577 1243 2631
<< m2 >>
rect 1197 2577 1243 2631
<< via1 >>
rect 1204 2584 1236 2624
<< m1 >>
rect 1197 2577 1243 2631
<< m2 >>
rect 1197 2577 1243 2631
<< via1 >>
rect 1204 2584 1236 2624
<< m1 >>
rect 685 1197 795 1251
<< m2 >>
rect 685 1197 795 1251
<< via1 >>
rect 692 1204 788 1244
<< m1 >>
rect 1261 1197 1371 1251
<< m2 >>
rect 1261 1197 1371 1251
<< via1 >>
rect 1268 1204 1364 1244
<< m1 >>
rect 1261 1197 1371 1251
<< m2 >>
rect 1261 1197 1371 1251
<< via1 >>
rect 1268 1204 1364 1244
<< m1 >>
rect 1453 517 1563 571
<< m2 >>
rect 1453 517 1563 571
<< via1 >>
rect 1460 524 1556 564
<< m1 >>
rect 1453 917 1563 971
<< m2 >>
rect 1453 917 1563 971
<< via1 >>
rect 1460 924 1556 964
<< m1 >>
rect 1197 2977 1243 3031
<< m2 >>
rect 1197 2977 1243 3031
<< via1 >>
rect 1204 2984 1236 3024
<< m1 >>
rect 1197 2977 1243 3031
<< m2 >>
rect 1197 2977 1243 3031
<< via1 >>
rect 1204 2984 1236 3024
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 1709 2417 1819 2471
<< m2 >>
rect 1709 2417 1819 2471
<< via1 >>
rect 1716 2424 1812 2464
<< m1 >>
rect 1709 2417 1819 2471
<< m2 >>
rect 1709 2417 1819 2471
<< m3 >>
rect 1709 2417 1819 2471
<< via2 >>
rect 1716 2424 1812 2464
<< via1 >>
rect 1716 2424 1812 2464
<< m1 >>
rect 877 3217 987 3271
<< m2 >>
rect 877 3217 987 3271
<< via1 >>
rect 884 3224 980 3264
<< m1 >>
rect 621 1477 667 1531
<< m2 >>
rect 621 1477 667 1531
<< via1 >>
rect 628 1484 660 1524
<< m1 >>
rect 621 1477 667 1531
<< m2 >>
rect 621 1477 667 1531
<< via1 >>
rect 628 1484 660 1524
<< m1 >>
rect 1197 1477 1243 1531
<< m2 >>
rect 1197 1477 1243 1531
<< via1 >>
rect 1204 1484 1236 1524
use COMP2 U1_COMP2 
transform 1 0 2298 0 1 0
box 0 0 1786 4158
use COMP3 U2_COMP3 
transform 1 0 4084 0 1 0
box 0 0 1786 4158
<< labels >>
flabel locali s 100 3958 2148 4008 0 FreeSans 400 0 0 0 VSS
port 4 nsew signal bidirectional
flabel locali s 0 4058 2248 4108 0 FreeSans 400 0 0 0 VDD
port 5 nsew signal bidirectional
flabel m1 s 628 1084 660 1124 0 FreeSans 400 0 0 0 VIP
port 6 nsew signal bidirectional
flabel m1 s 1204 1084 1236 1124 0 FreeSans 400 0 0 0 VIN
port 7 nsew signal bidirectional
flabel m2 s 930 2825 1521 2855 0 FreeSans 400 0 0 0 VO
port 8 nsew signal bidirectional
flabel m2 s 642 683 1218 713 0 FreeSans 400 0 0 0 I_BIAS
port 9 nsew signal bidirectional
<< properties >>
<< end >>
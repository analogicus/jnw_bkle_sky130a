magic
tech sky130A
magscale 1 1
timestamp 1748586004
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0  mirror1_MP2 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 504
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  mirror1_MP2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 264
box 0 0 576 240
use JNWATR_PCH_4C5F0  mirror1_MP1 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  mirror1_MP1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWATR_PCH_4C5F0  mirror1_MP3 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 2904
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mirror1_MP3_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 3304
box 0 0 576 240
use JNWATR_PCH_4C5F0  mirror3_MP4<9> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 904
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<8> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 904
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<7> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 2504
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<6> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 2504
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<5> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<4> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<3> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<2> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<1> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 1304
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP4<0> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 1304
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror3_MP5 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 2904
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mirror3_MP5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 3304
box 0 0 576 240
use JNWATR_NCH_4C5F0  None_MN1<9> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 4104
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  None_MN1<9>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 3864
box 0 0 576 240
use JNWATR_NCH_4C5F0  None_MN1<8> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 4104
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  None_MN1<8>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 3864
box 0 0 576 240
use JNWATR_NCH_4C5F0  None_MN1<7> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 5704
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN1<6> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 5704
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN1<5> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 5304
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN1<4> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 5304
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN1<3> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 6104
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  None_MN1<3>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 6504
box 0 0 576 240
use JNWATR_NCH_4C5F0  None_MN1<2> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 6104
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  None_MN1<2>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 6504
box 0 0 576 240
use JNWATR_NCH_4C5F0  None_MN1<1> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 4504
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN1<0> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 4504
box 0 0 576 400
use JNWATR_NCH_4C5F0  None_MN2 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 4904
box 0 0 576 400
use AALMISC_PNP_W3p40L3p40  diode_QP1 ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 6904
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<0> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 970 0 1 6904
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<1> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 9064
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<2> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 970 0 1 9064
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<3> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 8344
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<4> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 970 0 1 8344
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<5> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 7624
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<6> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 970 0 1 7624
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40  diode_QP2<7> ../AAL_MISC_SKY130A
timestamp 1748586004
transform 1 0 970 0 1 9784
box 0 0 670 670
use JNWATR_NCH_4C5F0  None_MN99 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 4904
box 0 0 576 400
<< m2 >>
rect 821 3085 964 3115
<< m3 >>
rect 821 685 851 3115
<< m2 >>
rect 821 685 979 715
<< m2 >>
rect 388 685 979 715
<< m2 >>
rect 814 3078 858 3122
<< m3 >>
rect 814 3078 858 3122
<< via2 >>
rect 821 3085 851 3115
<< m2 >>
rect 814 678 858 722
<< m3 >>
rect 814 678 858 722
<< via2 >>
rect 821 685 851 715
<< m2 >>
rect 1252 523 1411 553
<< m3 >>
rect 1381 523 1411 7129
<< m2 >>
rect 517 7099 1411 7129
<< m3 >>
rect 517 7099 547 7242
<< m2 >>
rect 1374 516 1418 560
<< m3 >>
rect 1374 516 1418 560
<< via2 >>
rect 1381 523 1411 553
<< m2 >>
rect 1374 7092 1418 7136
<< m3 >>
rect 1374 7092 1418 7136
<< via2 >>
rect 1381 7099 1411 7129
<< m2 >>
rect 510 7092 554 7136
<< m3 >>
rect 510 7092 554 7136
<< via2 >>
rect 517 7099 547 7129
<< m2 >>
rect 245 4288 388 4318
<< m3 >>
rect 245 4288 275 4718
<< m2 >>
rect 245 4688 403 4718
<< m2 >>
rect 245 4688 403 4718
<< m3 >>
rect 245 4688 275 5118
<< m2 >>
rect 245 5088 403 5118
<< m2 >>
rect 245 5088 403 5118
<< m3 >>
rect 245 5088 275 5518
<< m2 >>
rect 245 5488 403 5518
<< m2 >>
rect 245 5488 403 5518
<< m3 >>
rect 245 5488 275 5918
<< m2 >>
rect 245 5888 403 5918
<< m2 >>
rect 245 5888 403 5918
<< m3 >>
rect 245 5888 275 6318
<< m2 >>
rect 245 6288 403 6318
<< m2 >>
rect 373 6288 979 6318
<< m2 >>
rect 821 6288 979 6318
<< m3 >>
rect 821 5888 851 6318
<< m2 >>
rect 821 5888 979 5918
<< m2 >>
rect 821 5888 979 5918
<< m3 >>
rect 821 5488 851 5918
<< m2 >>
rect 821 5488 979 5518
<< m2 >>
rect 821 5488 979 5518
<< m3 >>
rect 821 4688 851 5518
<< m2 >>
rect 821 4688 979 4718
<< m2 >>
rect 821 4688 979 4718
<< m3 >>
rect 821 4288 851 4718
<< m2 >>
rect 821 4288 979 4318
<< m3 >>
rect 949 3296 979 4318
<< m2 >>
rect 949 3296 1267 3326
<< m3 >>
rect 1237 2943 1267 3326
<< m2 >>
rect 238 4281 282 4325
<< m3 >>
rect 238 4281 282 4325
<< via2 >>
rect 245 4288 275 4318
<< m2 >>
rect 238 4681 282 4725
<< m3 >>
rect 238 4681 282 4725
<< via2 >>
rect 245 4688 275 4718
<< m2 >>
rect 238 4681 282 4725
<< m3 >>
rect 238 4681 282 4725
<< via2 >>
rect 245 4688 275 4718
<< m2 >>
rect 238 5081 282 5125
<< m3 >>
rect 238 5081 282 5125
<< via2 >>
rect 245 5088 275 5118
<< m2 >>
rect 238 5081 282 5125
<< m3 >>
rect 238 5081 282 5125
<< via2 >>
rect 245 5088 275 5118
<< m2 >>
rect 238 5481 282 5525
<< m3 >>
rect 238 5481 282 5525
<< via2 >>
rect 245 5488 275 5518
<< m2 >>
rect 238 5481 282 5525
<< m3 >>
rect 238 5481 282 5525
<< via2 >>
rect 245 5488 275 5518
<< m2 >>
rect 238 5881 282 5925
<< m3 >>
rect 238 5881 282 5925
<< via2 >>
rect 245 5888 275 5918
<< m2 >>
rect 238 5881 282 5925
<< m3 >>
rect 238 5881 282 5925
<< via2 >>
rect 245 5888 275 5918
<< m2 >>
rect 238 6281 282 6325
<< m3 >>
rect 238 6281 282 6325
<< via2 >>
rect 245 6288 275 6318
<< m2 >>
rect 814 6281 858 6325
<< m3 >>
rect 814 6281 858 6325
<< via2 >>
rect 821 6288 851 6318
<< m2 >>
rect 814 5881 858 5925
<< m3 >>
rect 814 5881 858 5925
<< via2 >>
rect 821 5888 851 5918
<< m2 >>
rect 814 5881 858 5925
<< m3 >>
rect 814 5881 858 5925
<< via2 >>
rect 821 5888 851 5918
<< m2 >>
rect 814 5481 858 5525
<< m3 >>
rect 814 5481 858 5525
<< via2 >>
rect 821 5488 851 5518
<< m2 >>
rect 814 5481 858 5525
<< m3 >>
rect 814 5481 858 5525
<< via2 >>
rect 821 5488 851 5518
<< m2 >>
rect 814 4681 858 4725
<< m3 >>
rect 814 4681 858 4725
<< via2 >>
rect 821 4688 851 4718
<< m2 >>
rect 814 4681 858 4725
<< m3 >>
rect 814 4681 858 4725
<< via2 >>
rect 821 4688 851 4718
<< m2 >>
rect 814 4281 858 4325
<< m3 >>
rect 814 4281 858 4325
<< via2 >>
rect 821 4288 851 4318
<< m2 >>
rect 942 4281 986 4325
<< m3 >>
rect 942 4281 986 4325
<< via2 >>
rect 949 4288 979 4318
<< m2 >>
rect 942 3289 986 3333
<< m3 >>
rect 942 3289 986 3333
<< via2 >>
rect 949 3296 979 3326
<< m2 >>
rect 1230 3289 1274 3333
<< m3 >>
rect 1230 3289 1274 3333
<< via2 >>
rect 1237 3296 1267 3326
<< m2 >>
rect 149 4928 676 4958
<< m3 >>
rect 149 3088 179 4958
<< m2 >>
rect 149 3088 403 3118
<< m2 >>
rect 245 3088 403 3118
<< m3 >>
rect 245 2688 275 3118
<< m2 >>
rect 245 2688 403 2718
<< m2 >>
rect 245 2688 403 2718
<< m3 >>
rect 245 2288 275 2718
<< m2 >>
rect 245 2288 403 2318
<< m2 >>
rect 245 2288 403 2318
<< m3 >>
rect 245 1888 275 2318
<< m2 >>
rect 245 1888 403 1918
<< m2 >>
rect 245 1888 403 1918
<< m3 >>
rect 245 1488 275 1918
<< m2 >>
rect 245 1488 403 1518
<< m2 >>
rect 245 1488 403 1518
<< m3 >>
rect 245 1088 275 1518
<< m2 >>
rect 245 1088 403 1118
<< m2 >>
rect 373 1088 979 1118
<< m2 >>
rect 725 1088 979 1118
<< m3 >>
rect 725 1088 755 1246
<< m2 >>
rect 725 1216 947 1246
<< m3 >>
rect 917 1216 947 1390
<< m2 >>
rect 917 1360 1107 1390
<< m3 >>
rect 1077 1360 1107 1518
<< m2 >>
rect 949 1488 1107 1518
<< m2 >>
rect 725 1488 979 1518
<< m3 >>
rect 725 1488 755 1646
<< m2 >>
rect 725 1616 947 1646
<< m3 >>
rect 917 1616 947 1790
<< m2 >>
rect 917 1760 1107 1790
<< m3 >>
rect 1077 1760 1107 1918
<< m2 >>
rect 949 1888 1107 1918
<< m2 >>
rect 725 1888 979 1918
<< m3 >>
rect 725 1888 755 2046
<< m2 >>
rect 725 2016 947 2046
<< m3 >>
rect 917 2016 947 2190
<< m2 >>
rect 917 2160 1107 2190
<< m3 >>
rect 1077 2160 1107 2318
<< m2 >>
rect 949 2288 1107 2318
<< m2 >>
rect 725 2288 979 2318
<< m3 >>
rect 725 2288 755 2446
<< m2 >>
rect 725 2416 947 2446
<< m3 >>
rect 917 2416 947 2590
<< m2 >>
rect 917 2560 1107 2590
<< m3 >>
rect 1077 2560 1107 2718
<< m2 >>
rect 964 2688 1107 2718
<< m2 >>
rect 142 4921 186 4965
<< m3 >>
rect 142 4921 186 4965
<< via2 >>
rect 149 4928 179 4958
<< m2 >>
rect 142 3081 186 3125
<< m3 >>
rect 142 3081 186 3125
<< via2 >>
rect 149 3088 179 3118
<< m2 >>
rect 238 3081 282 3125
<< m3 >>
rect 238 3081 282 3125
<< via2 >>
rect 245 3088 275 3118
<< m2 >>
rect 238 2681 282 2725
<< m3 >>
rect 238 2681 282 2725
<< via2 >>
rect 245 2688 275 2718
<< m2 >>
rect 238 2681 282 2725
<< m3 >>
rect 238 2681 282 2725
<< via2 >>
rect 245 2688 275 2718
<< m2 >>
rect 238 2281 282 2325
<< m3 >>
rect 238 2281 282 2325
<< via2 >>
rect 245 2288 275 2318
<< m2 >>
rect 238 2281 282 2325
<< m3 >>
rect 238 2281 282 2325
<< via2 >>
rect 245 2288 275 2318
<< m2 >>
rect 238 1881 282 1925
<< m3 >>
rect 238 1881 282 1925
<< via2 >>
rect 245 1888 275 1918
<< m2 >>
rect 238 1881 282 1925
<< m3 >>
rect 238 1881 282 1925
<< via2 >>
rect 245 1888 275 1918
<< m2 >>
rect 238 1481 282 1525
<< m3 >>
rect 238 1481 282 1525
<< via2 >>
rect 245 1488 275 1518
<< m2 >>
rect 238 1481 282 1525
<< m3 >>
rect 238 1481 282 1525
<< via2 >>
rect 245 1488 275 1518
<< m2 >>
rect 238 1081 282 1125
<< m3 >>
rect 238 1081 282 1125
<< via2 >>
rect 245 1088 275 1118
<< m2 >>
rect 718 1081 762 1125
<< m3 >>
rect 718 1081 762 1125
<< via2 >>
rect 725 1088 755 1118
<< m2 >>
rect 718 1209 762 1253
<< m3 >>
rect 718 1209 762 1253
<< via2 >>
rect 725 1216 755 1246
<< m2 >>
rect 910 1209 954 1253
<< m3 >>
rect 910 1209 954 1253
<< via2 >>
rect 917 1216 947 1246
<< m2 >>
rect 910 1353 954 1397
<< m3 >>
rect 910 1353 954 1397
<< via2 >>
rect 917 1360 947 1390
<< m2 >>
rect 1070 1353 1114 1397
<< m3 >>
rect 1070 1353 1114 1397
<< via2 >>
rect 1077 1360 1107 1390
<< m2 >>
rect 1070 1481 1114 1525
<< m3 >>
rect 1070 1481 1114 1525
<< via2 >>
rect 1077 1488 1107 1518
<< m2 >>
rect 718 1481 762 1525
<< m3 >>
rect 718 1481 762 1525
<< via2 >>
rect 725 1488 755 1518
<< m2 >>
rect 718 1609 762 1653
<< m3 >>
rect 718 1609 762 1653
<< via2 >>
rect 725 1616 755 1646
<< m2 >>
rect 910 1609 954 1653
<< m3 >>
rect 910 1609 954 1653
<< via2 >>
rect 917 1616 947 1646
<< m2 >>
rect 910 1753 954 1797
<< m3 >>
rect 910 1753 954 1797
<< via2 >>
rect 917 1760 947 1790
<< m2 >>
rect 1070 1753 1114 1797
<< m3 >>
rect 1070 1753 1114 1797
<< via2 >>
rect 1077 1760 1107 1790
<< m2 >>
rect 1070 1881 1114 1925
<< m3 >>
rect 1070 1881 1114 1925
<< via2 >>
rect 1077 1888 1107 1918
<< m2 >>
rect 718 1881 762 1925
<< m3 >>
rect 718 1881 762 1925
<< via2 >>
rect 725 1888 755 1918
<< m2 >>
rect 718 2009 762 2053
<< m3 >>
rect 718 2009 762 2053
<< via2 >>
rect 725 2016 755 2046
<< m2 >>
rect 910 2009 954 2053
<< m3 >>
rect 910 2009 954 2053
<< via2 >>
rect 917 2016 947 2046
<< m2 >>
rect 910 2153 954 2197
<< m3 >>
rect 910 2153 954 2197
<< via2 >>
rect 917 2160 947 2190
<< m2 >>
rect 1070 2153 1114 2197
<< m3 >>
rect 1070 2153 1114 2197
<< via2 >>
rect 1077 2160 1107 2190
<< m2 >>
rect 1070 2281 1114 2325
<< m3 >>
rect 1070 2281 1114 2325
<< via2 >>
rect 1077 2288 1107 2318
<< m2 >>
rect 718 2281 762 2325
<< m3 >>
rect 718 2281 762 2325
<< via2 >>
rect 725 2288 755 2318
<< m2 >>
rect 718 2409 762 2453
<< m3 >>
rect 718 2409 762 2453
<< via2 >>
rect 725 2416 755 2446
<< m2 >>
rect 910 2409 954 2453
<< m3 >>
rect 910 2409 954 2453
<< via2 >>
rect 917 2416 947 2446
<< m2 >>
rect 910 2553 954 2597
<< m3 >>
rect 910 2553 954 2597
<< via2 >>
rect 917 2560 947 2590
<< m2 >>
rect 1070 2553 1114 2597
<< m3 >>
rect 1070 2553 1114 2597
<< via2 >>
rect 1077 2560 1107 2590
<< m2 >>
rect 1070 2681 1114 2725
<< m3 >>
rect 1070 2681 1114 2725
<< via2 >>
rect 1077 2688 1107 2718
<< m2 >>
rect 393 7947 536 7977
<< m3 >>
rect 393 7947 423 8697
<< m2 >>
rect 393 8667 551 8697
<< m2 >>
rect 393 8667 551 8697
<< m3 >>
rect 393 8667 423 9417
<< m2 >>
rect 393 9387 551 9417
<< m2 >>
rect 521 9387 1191 9417
<< m3 >>
rect 1161 9387 1191 10137
<< m2 >>
rect 1161 10107 1319 10137
<< m2 >>
rect 1289 10107 1447 10137
<< m3 >>
rect 1417 9387 1447 10137
<< m2 >>
rect 1289 9387 1447 9417
<< m2 >>
rect 1289 9387 1447 9417
<< m3 >>
rect 1417 8667 1447 9417
<< m2 >>
rect 1289 8667 1447 8697
<< m2 >>
rect 1289 8667 1447 8697
<< m3 >>
rect 1417 7947 1447 8697
<< m2 >>
rect 1289 7947 1447 7977
<< m2 >>
rect 1161 7947 1319 7977
<< m3 >>
rect 1161 7227 1191 7977
<< m2 >>
rect 1161 7227 1304 7257
<< m2 >>
rect 386 7940 430 7984
<< m3 >>
rect 386 7940 430 7984
<< via2 >>
rect 393 7947 423 7977
<< m2 >>
rect 386 8660 430 8704
<< m3 >>
rect 386 8660 430 8704
<< via2 >>
rect 393 8667 423 8697
<< m2 >>
rect 386 8660 430 8704
<< m3 >>
rect 386 8660 430 8704
<< via2 >>
rect 393 8667 423 8697
<< m2 >>
rect 386 9380 430 9424
<< m3 >>
rect 386 9380 430 9424
<< via2 >>
rect 393 9387 423 9417
<< m2 >>
rect 1154 9380 1198 9424
<< m3 >>
rect 1154 9380 1198 9424
<< via2 >>
rect 1161 9387 1191 9417
<< m2 >>
rect 1154 10100 1198 10144
<< m3 >>
rect 1154 10100 1198 10144
<< via2 >>
rect 1161 10107 1191 10137
<< m2 >>
rect 1410 10100 1454 10144
<< m3 >>
rect 1410 10100 1454 10144
<< via2 >>
rect 1417 10107 1447 10137
<< m2 >>
rect 1410 9380 1454 9424
<< m3 >>
rect 1410 9380 1454 9424
<< via2 >>
rect 1417 9387 1447 9417
<< m2 >>
rect 1410 9380 1454 9424
<< m3 >>
rect 1410 9380 1454 9424
<< via2 >>
rect 1417 9387 1447 9417
<< m2 >>
rect 1410 8660 1454 8704
<< m3 >>
rect 1410 8660 1454 8704
<< via2 >>
rect 1417 8667 1447 8697
<< m2 >>
rect 1410 8660 1454 8704
<< m3 >>
rect 1410 8660 1454 8704
<< via2 >>
rect 1417 8667 1447 8697
<< m2 >>
rect 1410 7940 1454 7984
<< m3 >>
rect 1410 7940 1454 7984
<< via2 >>
rect 1417 7947 1447 7977
<< m2 >>
rect 1154 7940 1198 7984
<< m3 >>
rect 1154 7940 1198 7984
<< via2 >>
rect 1161 7947 1191 7977
<< m2 >>
rect 1154 7220 1198 7264
<< m3 >>
rect 1154 7220 1198 7264
<< via2 >>
rect 1161 7227 1191 7257
<< locali >>
rect 100 10504 1740 10554
<< locali >>
rect 100 100 1740 150
<< m1 >>
rect 100 150 150 10504
<< m1 >>
rect 1690 150 1740 10504
<< locali >>
rect 93 10497 157 10561
<< m1 >>
rect 93 10497 157 10561
<< viali >>
rect 100 10504 150 10554
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1683 10497 1747 10561
<< m1 >>
rect 1683 10497 1747 10561
<< viali >>
rect 1690 10504 1740 10554
<< locali >>
rect 1683 93 1747 157
<< m1 >>
rect 1683 93 1747 157
<< viali >>
rect 1690 100 1740 150
<< locali >>
rect 0 10604 1840 10654
<< locali >>
rect 0 0 1840 50
<< m1 >>
rect 0 50 50 10604
<< m1 >>
rect 1790 50 1840 10604
<< locali >>
rect -7 10597 57 10661
<< m1 >>
rect -7 10597 57 10661
<< viali >>
rect 0 10604 50 10654
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1783 10597 1847 10661
<< m1 >>
rect 1783 10597 1847 10661
<< viali >>
rect 1790 10604 1840 10654
<< locali >>
rect 1783 -7 1847 57
<< m1 >>
rect 1783 -7 1847 57
<< viali >>
rect 1790 0 1840 50
<< locali >>
rect 244 804 532 844
<< locali >>
rect 820 804 1108 844
<< locali >>
rect 820 3204 1108 3244
<< locali >>
rect 820 1204 1108 1244
<< locali >>
rect 1204 1084 1364 1124
<< locali >>
rect 244 1204 532 1244
<< locali >>
rect 628 1084 788 1124
<< locali >>
rect 820 2804 1108 2844
<< locali >>
rect 1204 2684 1364 2724
<< locali >>
rect 244 2804 532 2844
<< locali >>
rect 628 2684 788 2724
<< locali >>
rect 820 2004 1108 2044
<< locali >>
rect 1204 1884 1364 1924
<< locali >>
rect 244 2004 532 2044
<< locali >>
rect 628 1884 788 1924
<< locali >>
rect 820 2404 1108 2444
<< locali >>
rect 1204 2284 1364 2324
<< locali >>
rect 244 2404 532 2444
<< locali >>
rect 628 2284 788 2324
<< locali >>
rect 244 1604 532 1644
<< locali >>
rect 628 1484 788 1524
<< locali >>
rect 820 1604 1108 1644
<< locali >>
rect 1204 1484 1364 1524
<< locali >>
rect 244 3204 532 3244
<< locali >>
rect 820 4404 1108 4444
<< locali >>
rect 1204 4284 1364 4324
<< locali >>
rect 244 4404 532 4444
<< locali >>
rect 628 4284 788 4324
<< locali >>
rect 244 6004 532 6044
<< locali >>
rect 628 5884 788 5924
<< locali >>
rect 820 6004 1108 6044
<< locali >>
rect 1204 5884 1364 5924
<< locali >>
rect 244 5604 532 5644
<< locali >>
rect 628 5484 788 5524
<< locali >>
rect 820 5604 1108 5644
<< locali >>
rect 1204 5484 1364 5524
<< locali >>
rect 244 6404 532 6444
<< locali >>
rect 628 6284 788 6324
<< locali >>
rect 820 6404 1108 6444
<< locali >>
rect 1204 6284 1364 6324
<< locali >>
rect 244 4804 532 4844
<< locali >>
rect 628 4684 788 4724
<< locali >>
rect 820 4804 1108 4844
<< locali >>
rect 1204 4684 1364 4724
<< locali >>
rect 244 5204 532 5244
<< locali >>
rect 820 5204 1108 5244
<< locali >>
rect 0 336 1840 432
<< locali >>
rect -7 329 57 439
<< m1 >>
rect -7 329 57 439
<< viali >>
rect 0 336 50 432
<< locali >>
rect 1783 329 1847 439
<< m1 >>
rect 1783 329 1847 439
<< viali >>
rect 1790 336 1840 432
<< locali >>
rect 0 3376 1840 3472
<< locali >>
rect -7 3369 57 3479
<< m1 >>
rect -7 3369 57 3479
<< viali >>
rect 0 3376 50 3472
<< locali >>
rect 1783 3369 1847 3479
<< m1 >>
rect 1783 3369 1847 3479
<< viali >>
rect 1790 3376 1840 3472
<< locali >>
rect 100 3936 1740 4032
<< locali >>
rect 93 3929 157 4039
<< m1 >>
rect 93 3929 157 4039
<< viali >>
rect 100 3936 150 4032
<< locali >>
rect 1683 3929 1747 4039
<< m1 >>
rect 1683 3929 1747 4039
<< viali >>
rect 1690 3936 1740 4032
<< locali >>
rect 100 6576 1740 6672
<< locali >>
rect 93 6569 157 6679
<< m1 >>
rect 93 6569 157 6679
<< viali >>
rect 100 6576 150 6672
<< locali >>
rect 1683 6569 1747 6679
<< m1 >>
rect 1683 6569 1747 6679
<< viali >>
rect 1690 6576 1740 6672
<< locali >>
rect 510 7479 560 7512
<< locali >>
rect 1280 7479 1330 7512
<< locali >>
rect 510 9639 560 9672
<< locali >>
rect 1280 9639 1330 9672
<< locali >>
rect 510 8919 560 8952
<< locali >>
rect 1280 8919 1330 8952
<< locali >>
rect 510 8199 560 8232
<< locali >>
rect 1280 8199 1330 8232
<< locali >>
rect 1280 10359 1330 10392
<< locali >>
rect 100 7525 1740 7574
<< locali >>
rect 93 7518 157 7581
<< m1 >>
rect 93 7518 157 7581
<< viali >>
rect 100 7525 150 7574
<< locali >>
rect 1683 7518 1747 7581
<< m1 >>
rect 1683 7518 1747 7581
<< viali >>
rect 1690 7525 1740 7574
<< locali >>
rect 100 6904 1740 6953
<< locali >>
rect 93 6897 157 6960
<< m1 >>
rect 93 6897 157 6960
<< viali >>
rect 100 6904 150 6953
<< locali >>
rect 1683 6897 1747 6960
<< m1 >>
rect 1683 6897 1747 6960
<< viali >>
rect 1690 6904 1740 6953
<< locali >>
rect 100 9685 1740 9734
<< locali >>
rect 93 9678 157 9741
<< m1 >>
rect 93 9678 157 9741
<< viali >>
rect 100 9685 150 9734
<< locali >>
rect 1683 9678 1747 9741
<< m1 >>
rect 1683 9678 1747 9741
<< viali >>
rect 1690 9685 1740 9734
<< locali >>
rect 100 9064 1740 9113
<< locali >>
rect 93 9057 157 9120
<< m1 >>
rect 93 9057 157 9120
<< viali >>
rect 100 9064 150 9113
<< locali >>
rect 1683 9057 1747 9120
<< m1 >>
rect 1683 9057 1747 9120
<< viali >>
rect 1690 9064 1740 9113
<< locali >>
rect 100 8965 1740 9014
<< locali >>
rect 93 8958 157 9021
<< m1 >>
rect 93 8958 157 9021
<< viali >>
rect 100 8965 150 9014
<< locali >>
rect 1683 8958 1747 9021
<< m1 >>
rect 1683 8958 1747 9021
<< viali >>
rect 1690 8965 1740 9014
<< locali >>
rect 100 8344 1740 8393
<< locali >>
rect 93 8337 157 8400
<< m1 >>
rect 93 8337 157 8400
<< viali >>
rect 100 8344 150 8393
<< locali >>
rect 1683 8337 1747 8400
<< m1 >>
rect 1683 8337 1747 8400
<< viali >>
rect 1690 8344 1740 8393
<< locali >>
rect 100 8245 1740 8294
<< locali >>
rect 93 8238 157 8301
<< m1 >>
rect 93 8238 157 8301
<< viali >>
rect 100 8245 150 8294
<< locali >>
rect 1683 8238 1747 8301
<< m1 >>
rect 1683 8238 1747 8301
<< viali >>
rect 1690 8245 1740 8294
<< locali >>
rect 100 7624 1740 7673
<< locali >>
rect 93 7617 157 7680
<< m1 >>
rect 93 7617 157 7680
<< viali >>
rect 100 7624 150 7673
<< locali >>
rect 1683 7617 1747 7680
<< m1 >>
rect 1683 7617 1747 7680
<< viali >>
rect 1690 7624 1740 7673
<< locali >>
rect 100 10405 1740 10454
<< locali >>
rect 93 10398 157 10461
<< m1 >>
rect 93 10398 157 10461
<< viali >>
rect 100 10405 150 10454
<< locali >>
rect 1683 10398 1747 10461
<< m1 >>
rect 1683 10398 1747 10461
<< viali >>
rect 1690 10405 1740 10454
<< locali >>
rect 100 9784 1740 9833
<< locali >>
rect 93 9777 157 9840
<< m1 >>
rect 93 9777 157 9840
<< viali >>
rect 100 9784 150 9833
<< locali >>
rect 1683 9777 1747 9840
<< m1 >>
rect 1683 9777 1747 9840
<< viali >>
rect 1690 9784 1740 9833
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 3077 987 3131
<< m2 >>
rect 941 3077 987 3131
<< via1 >>
rect 948 3084 980 3124
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 483 7210 587 7276
<< m2 >>
rect 483 7210 587 7276
<< m3 >>
rect 483 7210 587 7276
<< via2 >>
rect 490 7217 580 7269
<< via1 >>
rect 490 7217 580 7269
<< m1 >>
rect 1197 2917 1307 2971
<< m2 >>
rect 1197 2917 1307 2971
<< m3 >>
rect 1197 2917 1307 2971
<< via2 >>
rect 1204 2924 1300 2964
<< via1 >>
rect 1204 2924 1300 2964
<< m1 >>
rect 941 4277 987 4331
<< m2 >>
rect 941 4277 987 4331
<< via1 >>
rect 948 4284 980 4324
<< m1 >>
rect 941 4277 987 4331
<< m2 >>
rect 941 4277 987 4331
<< m3 >>
rect 941 4277 987 4331
<< via2 >>
rect 948 4284 980 4324
<< via1 >>
rect 948 4284 980 4324
<< m1 >>
rect 365 4277 411 4331
<< m2 >>
rect 365 4277 411 4331
<< via1 >>
rect 372 4284 404 4324
<< m1 >>
rect 365 5877 411 5931
<< m2 >>
rect 365 5877 411 5931
<< via1 >>
rect 372 5884 404 5924
<< m1 >>
rect 365 5877 411 5931
<< m2 >>
rect 365 5877 411 5931
<< via1 >>
rect 372 5884 404 5924
<< m1 >>
rect 941 5877 987 5931
<< m2 >>
rect 941 5877 987 5931
<< via1 >>
rect 948 5884 980 5924
<< m1 >>
rect 941 5877 987 5931
<< m2 >>
rect 941 5877 987 5931
<< via1 >>
rect 948 5884 980 5924
<< m1 >>
rect 365 5477 411 5531
<< m2 >>
rect 365 5477 411 5531
<< via1 >>
rect 372 5484 404 5524
<< m1 >>
rect 365 5477 411 5531
<< m2 >>
rect 365 5477 411 5531
<< via1 >>
rect 372 5484 404 5524
<< m1 >>
rect 941 5477 987 5531
<< m2 >>
rect 941 5477 987 5531
<< via1 >>
rect 948 5484 980 5524
<< m1 >>
rect 941 5477 987 5531
<< m2 >>
rect 941 5477 987 5531
<< via1 >>
rect 948 5484 980 5524
<< m1 >>
rect 365 6277 411 6331
<< m2 >>
rect 365 6277 411 6331
<< via1 >>
rect 372 6284 404 6324
<< m1 >>
rect 365 6277 411 6331
<< m2 >>
rect 365 6277 411 6331
<< via1 >>
rect 372 6284 404 6324
<< m1 >>
rect 941 6277 987 6331
<< m2 >>
rect 941 6277 987 6331
<< via1 >>
rect 948 6284 980 6324
<< m1 >>
rect 941 6277 987 6331
<< m2 >>
rect 941 6277 987 6331
<< via1 >>
rect 948 6284 980 6324
<< m1 >>
rect 365 4677 411 4731
<< m2 >>
rect 365 4677 411 4731
<< via1 >>
rect 372 4684 404 4724
<< m1 >>
rect 365 4677 411 4731
<< m2 >>
rect 365 4677 411 4731
<< via1 >>
rect 372 4684 404 4724
<< m1 >>
rect 941 4677 987 4731
<< m2 >>
rect 941 4677 987 4731
<< via1 >>
rect 948 4684 980 4724
<< m1 >>
rect 941 4677 987 4731
<< m2 >>
rect 941 4677 987 4731
<< via1 >>
rect 948 4684 980 4724
<< m1 >>
rect 365 5077 411 5131
<< m2 >>
rect 365 5077 411 5131
<< via1 >>
rect 372 5084 404 5124
<< m1 >>
rect 365 5077 411 5131
<< m2 >>
rect 365 5077 411 5131
<< via1 >>
rect 372 5084 404 5124
<< m1 >>
rect 941 1077 987 1131
<< m2 >>
rect 941 1077 987 1131
<< via1 >>
rect 948 1084 980 1124
<< m1 >>
rect 941 1077 987 1131
<< m2 >>
rect 941 1077 987 1131
<< via1 >>
rect 948 1084 980 1124
<< m1 >>
rect 365 1077 411 1131
<< m2 >>
rect 365 1077 411 1131
<< via1 >>
rect 372 1084 404 1124
<< m1 >>
rect 365 1077 411 1131
<< m2 >>
rect 365 1077 411 1131
<< via1 >>
rect 372 1084 404 1124
<< m1 >>
rect 941 2677 987 2731
<< m2 >>
rect 941 2677 987 2731
<< via1 >>
rect 948 2684 980 2724
<< m1 >>
rect 365 2677 411 2731
<< m2 >>
rect 365 2677 411 2731
<< via1 >>
rect 372 2684 404 2724
<< m1 >>
rect 365 2677 411 2731
<< m2 >>
rect 365 2677 411 2731
<< via1 >>
rect 372 2684 404 2724
<< m1 >>
rect 941 1877 987 1931
<< m2 >>
rect 941 1877 987 1931
<< via1 >>
rect 948 1884 980 1924
<< m1 >>
rect 941 1877 987 1931
<< m2 >>
rect 941 1877 987 1931
<< via1 >>
rect 948 1884 980 1924
<< m1 >>
rect 365 1877 411 1931
<< m2 >>
rect 365 1877 411 1931
<< via1 >>
rect 372 1884 404 1924
<< m1 >>
rect 365 1877 411 1931
<< m2 >>
rect 365 1877 411 1931
<< via1 >>
rect 372 1884 404 1924
<< m1 >>
rect 941 2277 987 2331
<< m2 >>
rect 941 2277 987 2331
<< via1 >>
rect 948 2284 980 2324
<< m1 >>
rect 941 2277 987 2331
<< m2 >>
rect 941 2277 987 2331
<< via1 >>
rect 948 2284 980 2324
<< m1 >>
rect 365 2277 411 2331
<< m2 >>
rect 365 2277 411 2331
<< via1 >>
rect 372 2284 404 2324
<< m1 >>
rect 365 2277 411 2331
<< m2 >>
rect 365 2277 411 2331
<< via1 >>
rect 372 2284 404 2324
<< m1 >>
rect 365 1477 411 1531
<< m2 >>
rect 365 1477 411 1531
<< via1 >>
rect 372 1484 404 1524
<< m1 >>
rect 365 1477 411 1531
<< m2 >>
rect 365 1477 411 1531
<< via1 >>
rect 372 1484 404 1524
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 365 3077 411 3131
<< m2 >>
rect 365 3077 411 3131
<< via1 >>
rect 372 3084 404 3124
<< m1 >>
rect 365 3077 411 3131
<< m2 >>
rect 365 3077 411 3131
<< via1 >>
rect 372 3084 404 3124
<< m1 >>
rect 621 4917 731 4971
<< m2 >>
rect 621 4917 731 4971
<< via1 >>
rect 628 4924 724 4964
<< m1 >>
rect 1253 7210 1357 7276
<< m2 >>
rect 1253 7210 1357 7276
<< via1 >>
rect 1260 7217 1350 7269
<< m1 >>
rect 483 9370 587 9436
<< m2 >>
rect 483 9370 587 9436
<< via1 >>
rect 490 9377 580 9429
<< m1 >>
rect 483 9370 587 9436
<< m2 >>
rect 483 9370 587 9436
<< via1 >>
rect 490 9377 580 9429
<< m1 >>
rect 1253 9370 1357 9436
<< m2 >>
rect 1253 9370 1357 9436
<< via1 >>
rect 1260 9377 1350 9429
<< m1 >>
rect 1253 9370 1357 9436
<< m2 >>
rect 1253 9370 1357 9436
<< via1 >>
rect 1260 9377 1350 9429
<< m1 >>
rect 483 8650 587 8716
<< m2 >>
rect 483 8650 587 8716
<< via1 >>
rect 490 8657 580 8709
<< m1 >>
rect 483 8650 587 8716
<< m2 >>
rect 483 8650 587 8716
<< via1 >>
rect 490 8657 580 8709
<< m1 >>
rect 1253 8650 1357 8716
<< m2 >>
rect 1253 8650 1357 8716
<< via1 >>
rect 1260 8657 1350 8709
<< m1 >>
rect 1253 8650 1357 8716
<< m2 >>
rect 1253 8650 1357 8716
<< via1 >>
rect 1260 8657 1350 8709
<< m1 >>
rect 483 7930 587 7996
<< m2 >>
rect 483 7930 587 7996
<< via1 >>
rect 490 7937 580 7989
<< m1 >>
rect 1253 7930 1357 7996
<< m2 >>
rect 1253 7930 1357 7996
<< via1 >>
rect 1260 7937 1350 7989
<< m1 >>
rect 1253 7930 1357 7996
<< m2 >>
rect 1253 7930 1357 7996
<< via1 >>
rect 1260 7937 1350 7989
<< m1 >>
rect 1253 10090 1357 10156
<< m2 >>
rect 1253 10090 1357 10156
<< via1 >>
rect 1260 10097 1350 10149
<< m1 >>
rect 1253 10090 1357 10156
<< m2 >>
rect 1253 10090 1357 10156
<< via1 >>
rect 1260 10097 1350 10149
use OTA U1_OTA 
transform 1 0 1890 0 1 0
box 0 0 2686 9614
use JNW_BKLE_GR06_res U2_JNW_BKLE_GR06_res 
transform 1 0 4576 0 1 0
box 0 0 1390 6952
<< labels >>
flabel locali s 0 10604 1840 10654 0 FreeSans 400 0 0 0 VDD
port 35 nsew signal bidirectional
flabel locali s 100 10504 1740 10554 0 FreeSans 400 0 0 0 VSS
port 36 nsew signal bidirectional
flabel m1 s 628 2924 724 2964 0 FreeSans 400 0 0 0 OUT
port 37 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744575209
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 2600
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 2360
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 2600
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 2360
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 360
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 360
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1800
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 1800
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3800
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 3400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 3800
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3000
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1000
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 976 0 1 1000
box 0 0 576 400
<< locali >>
rect 150 4150 1802 4250
<< locali >>
rect 150 150 1802 250
<< m1 >>
rect 150 250 250 4150
<< m1 >>
rect 1702 250 1802 4150
<< locali >>
rect 143 4143 257 4257
<< m1 >>
rect 143 4143 257 4257
<< viali >>
rect 150 4150 250 4250
<< locali >>
rect 143 143 257 257
<< m1 >>
rect 143 143 257 257
<< viali >>
rect 150 150 250 250
<< locali >>
rect 1695 4143 1809 4257
<< m1 >>
rect 1695 4143 1809 4257
<< viali >>
rect 1702 4150 1802 4250
<< locali >>
rect 1695 143 1809 257
<< m1 >>
rect 1695 143 1809 257
<< viali >>
rect 1702 150 1802 250
<< locali >>
rect 0 4300 1952 4400
<< locali >>
rect 0 0 1952 100
<< m1 >>
rect 0 100 100 4300
<< m1 >>
rect 1852 100 1952 4300
<< locali >>
rect -7 4293 107 4407
<< m1 >>
rect -7 4293 107 4407
<< viali >>
rect 0 4300 100 4400
<< locali >>
rect -7 -7 107 107
<< m1 >>
rect -7 -7 107 107
<< viali >>
rect 0 0 100 100
<< locali >>
rect 1845 4293 1959 4407
<< m1 >>
rect 1845 4293 1959 4407
<< viali >>
rect 1852 4300 1952 4400
<< locali >>
rect 1845 -7 1959 107
<< m1 >>
rect 1845 -7 1959 107
<< viali >>
rect 1852 0 1952 100
<< locali >>
rect 352 900 640 940
<< locali >>
rect 736 780 896 820
<< locali >>
rect 928 900 1216 940
<< locali >>
rect 352 1700 640 1740
<< locali >>
rect 928 1700 1216 1740
<< locali >>
rect 1312 1580 1472 1620
<< locali >>
rect 352 3700 640 3740
<< locali >>
rect 928 3700 1216 3740
<< locali >>
rect 1312 3580 1472 3620
<< locali >>
rect 352 3300 640 3340
<< locali >>
rect 736 3180 896 3220
<< locali >>
rect 928 3300 1216 3340
<< locali >>
rect 352 1300 640 1340
<< locali >>
rect 928 1300 1216 1340
<< locali >>
rect 0 2432 1952 2528
<< locali >>
rect -7 2425 107 2535
<< m1 >>
rect -7 2425 107 2535
<< viali >>
rect 0 2432 100 2528
<< locali >>
rect 1845 2425 1959 2535
<< m1 >>
rect 1845 2425 1959 2535
<< viali >>
rect 1852 2432 1952 2528
<< locali >>
rect 150 432 1802 528
<< locali >>
rect 143 425 257 535
<< m1 >>
rect 143 425 257 535
<< viali >>
rect 150 432 250 528
<< locali >>
rect 1695 425 1809 535
<< m1 >>
rect 1695 425 1809 535
<< viali >>
rect 1702 432 1802 528
<< locali >>
rect 150 1872 1802 1968
<< locali >>
rect 143 1865 257 1975
<< m1 >>
rect 143 1865 257 1975
<< viali >>
rect 150 1872 250 1968
<< locali >>
rect 1695 1865 1809 1975
<< m1 >>
rect 1695 1865 1809 1975
<< viali >>
rect 1702 1872 1802 1968
<< locali >>
rect 0 3872 1952 3968
<< locali >>
rect -7 3865 107 3975
<< m1 >>
rect -7 3865 107 3975
<< viali >>
rect 0 3872 100 3968
<< locali >>
rect 1845 3865 1959 3975
<< m1 >>
rect 1845 3865 1959 3975
<< viali >>
rect 1852 3872 1952 3968
<< labels >>
flabel locali s 0 4300 1952 4400 0 FreeSans 400 0 0 0 VSS
port 44 nsew signal bidirectional
flabel locali s 150 4150 1802 4250 0 FreeSans 400 0 0 0 VDD
port 45 nsew signal bidirectional
<< properties >>
<< end >>
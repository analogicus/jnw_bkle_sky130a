magic
tech sky130A
magscale 1 1
timestamp 1729517738
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 x1 ../JNW_ATR_SKY130A
transform 0 1 2500 -1 0 1500
box 0 0 832 400
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform 0 1 4000 -1 0 1500
box 0 0 512 400
use JNWTR_RES2 x3 ../JNW_TR_SKY130A
transform 0 1 5500 -1 0 1500
box 0 0 324 1320
use JNWATR_NCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 0 1 7000 -1 0 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x3 ../JNW_ATR_SKY130A
transform 0 1 8500 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x7 ../JNW_ATR_SKY130A
transform 0 1 10000 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x9 ../JNW_ATR_SKY130A
transform 0 1 11500 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x8 ../JNW_ATR_SKY130A
transform 0 1 13000 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x5 ../JNW_ATR_SKY130A
transform 0 1 14500 -1 0 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform 0 1 16000 -1 0 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 0 1 17500 -1 0 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x10 ../JNW_ATR_SKY130A
transform 0 1 19000 -1 0 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x11 ../JNW_ATR_SKY130A
transform 0 1 20500 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x12 ../JNW_ATR_SKY130A
transform 0 1 22000 -1 0 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x13 ../JNW_ATR_SKY130A
transform 0 1 23500 -1 0 1500
box 0 0 576 400
<< labels >>
<< properties >>
<< end >>
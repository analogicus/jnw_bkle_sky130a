magic
tech sky130A
magscale 1 1
timestamp 1746712773
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2804
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2804
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1604
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1364
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1604
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1364
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 3604
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 3604
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 264
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 7504
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 5724
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 3954
box 0 0 2236 1720
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 941 2977 987 3031
<< m2 >>
rect 941 2977 987 3031
<< via1 >>
rect 948 2984 980 3024
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< m3 >>
rect 365 2577 411 2631
<< via2 >>
rect 372 2584 404 2624
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< m3 >>
rect 941 2577 987 2631
<< via2 >>
rect 948 2584 980 2624
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 365 1777 411 1831
<< m2 >>
rect 365 1777 411 1831
<< via1 >>
rect 372 1784 404 1824
<< m1 >>
rect 941 1777 987 1831
<< m2 >>
rect 941 1777 987 1831
<< via1 >>
rect 948 1784 980 1824
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< m3 >>
rect 365 2177 411 2231
<< via2 >>
rect 372 2184 404 2224
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< m3 >>
rect 941 2177 987 2231
<< via2 >>
rect 948 2184 980 2224
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< m3 >>
rect 621 1617 731 1671
<< via2 >>
rect 628 1624 724 1664
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< m3 >>
rect 621 1617 731 1671
<< via2 >>
rect 628 1624 724 1664
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< m3 >>
rect 621 1617 731 1671
<< via2 >>
rect 628 1624 724 1664
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 1197 1617 1307 1671
<< m2 >>
rect 1197 1617 1307 1671
<< m3 >>
rect 1197 1617 1307 1671
<< via2 >>
rect 1204 1624 1300 1664
<< via1 >>
rect 1204 1624 1300 1664
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< m3 >>
rect 621 2017 731 2071
<< via2 >>
rect 628 2024 724 2064
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< m3 >>
rect 621 2017 731 2071
<< via2 >>
rect 628 2024 724 2064
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< m3 >>
rect 1197 2017 1307 2071
<< via2 >>
rect 1204 2024 1300 2064
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< m3 >>
rect 1197 2017 1307 2071
<< via2 >>
rect 1204 2024 1300 2064
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 621 517 731 571
<< m2 >>
rect 621 517 731 571
<< m3 >>
rect 621 517 731 571
<< via2 >>
rect 628 524 724 564
<< via1 >>
rect 628 524 724 564
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< m3 >>
rect 621 2817 731 2871
<< via2 >>
rect 628 2824 724 2864
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< m3 >>
rect 621 2817 731 2871
<< via2 >>
rect 628 2824 724 2864
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< m3 >>
rect 1197 2817 1307 2871
<< via2 >>
rect 1204 2824 1300 2864
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< m3 >>
rect 1197 2817 1307 2871
<< via2 >>
rect 1204 2824 1300 2864
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 621 2417 731 2471
<< m2 >>
rect 621 2417 731 2471
<< m3 >>
rect 621 2417 731 2471
<< via2 >>
rect 628 2424 724 2464
<< via1 >>
rect 628 2424 724 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< m3 >>
rect 1197 2417 1307 2471
<< via2 >>
rect 1204 2424 1300 2464
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< m3 >>
rect 1197 2417 1307 2471
<< via2 >>
rect 1204 2424 1300 2464
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< m3 >>
rect 941 677 987 731
<< via2 >>
rect 948 684 980 724
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< m3 >>
rect 941 677 987 731
<< via2 >>
rect 948 684 980 724
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< m3 >>
rect 1197 517 1307 571
<< via2 >>
rect 1204 524 1300 564
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< m3 >>
rect 429 3097 539 3151
<< via2 >>
rect 436 3104 532 3144
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 1005 3097 1115 3151
<< m2 >>
rect 1005 3097 1115 3151
<< via1 >>
rect 1012 3104 1108 3144
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< m3 >>
rect 429 2697 539 2751
<< via2 >>
rect 436 2704 532 2744
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< m3 >>
rect 1005 2697 1115 2751
<< via2 >>
rect 1012 2704 1108 2744
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< m3 >>
rect 429 1897 539 1951
<< via2 >>
rect 436 1904 532 1944
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< m3 >>
rect 1005 1897 1115 1951
<< via2 >>
rect 1012 1904 1108 1944
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< m3 >>
rect 429 2297 539 2351
<< via2 >>
rect 436 2304 532 2344
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< m3 >>
rect 1005 2297 1115 2351
<< via2 >>
rect 1012 2304 1108 2344
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1197 3217 1307 3271
<< m2 >>
rect 1197 3217 1307 3271
<< via1 >>
rect 1204 3224 1300 3264
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< m3 >>
rect 941 3377 987 3431
<< via2 >>
rect 948 3384 980 3424
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< m3 >>
rect 941 3377 987 3431
<< via2 >>
rect 948 3384 980 3424
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 621 3217 731 3271
<< m2 >>
rect 621 3217 731 3271
<< via1 >>
rect 628 3224 724 3264
<< locali >>
rect 2103 8957 2261 9091
<< m1 >>
rect 2103 8957 2261 9091
<< m2 >>
rect 2103 8957 2261 9091
<< via1 >>
rect 2110 8964 2254 9084
<< viali >>
rect 2110 8964 2254 9084
<< locali >>
rect 375 8957 533 9091
<< m1 >>
rect 375 8957 533 9091
<< m2 >>
rect 375 8957 533 9091
<< m3 >>
rect 375 8957 533 9091
<< via2 >>
rect 382 8964 526 9084
<< via1 >>
rect 382 8964 526 9084
<< viali >>
rect 382 8964 526 9084
<< locali >>
rect 2103 7177 2261 7311
<< m1 >>
rect 2103 7177 2261 7311
<< m2 >>
rect 2103 7177 2261 7311
<< m3 >>
rect 2103 7177 2261 7311
<< via2 >>
rect 2110 7184 2254 7304
<< via1 >>
rect 2110 7184 2254 7304
<< viali >>
rect 2110 7184 2254 7304
<< locali >>
rect 375 7177 533 7311
<< m1 >>
rect 375 7177 533 7311
<< m2 >>
rect 375 7177 533 7311
<< m3 >>
rect 375 7177 533 7311
<< via2 >>
rect 382 7184 526 7304
<< via1 >>
rect 382 7184 526 7304
<< viali >>
rect 382 7184 526 7304
<< locali >>
rect 2103 5407 2261 5541
<< m1 >>
rect 2103 5407 2261 5541
<< m2 >>
rect 2103 5407 2261 5541
<< m3 >>
rect 2103 5407 2261 5541
<< via2 >>
rect 2110 5414 2254 5534
<< via1 >>
rect 2110 5414 2254 5534
<< viali >>
rect 2110 5414 2254 5534
<< m2 >>
rect 819 2987 962 3017
<< m3 >>
rect 819 2587 849 3017
<< m2 >>
rect 819 2587 977 2617
<< m3 >>
rect 947 2587 977 2617
<< m2 >>
rect 371 2587 977 2617
<< m3 >>
rect 371 2587 401 2617
<< m2 >>
rect 243 2587 401 2617
<< m3 >>
rect 243 2587 273 3017
<< m2 >>
rect 243 2987 386 3017
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 941 2977 987 3031
<< m2 >>
rect 941 2977 987 3031
<< via1 >>
rect 948 2984 980 3024
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m2 >>
rect 812 2980 856 3024
<< m3 >>
rect 812 2980 856 3024
<< via2 >>
rect 819 2987 849 3017
<< m2 >>
rect 812 2580 856 2624
<< m3 >>
rect 812 2580 856 2624
<< via2 >>
rect 819 2587 849 2617
<< m2 >>
rect 940 2580 984 2624
<< m3 >>
rect 940 2580 984 2624
<< via2 >>
rect 947 2587 977 2617
<< m2 >>
rect 940 2580 984 2624
<< m3 >>
rect 940 2580 984 2624
<< via2 >>
rect 947 2587 977 2617
<< m2 >>
rect 364 2580 408 2624
<< m3 >>
rect 364 2580 408 2624
<< via2 >>
rect 371 2587 401 2617
<< m2 >>
rect 364 2580 408 2624
<< m3 >>
rect 364 2580 408 2624
<< via2 >>
rect 371 2587 401 2617
<< m2 >>
rect 236 2580 280 2624
<< m3 >>
rect 236 2580 280 2624
<< via2 >>
rect 243 2587 273 2617
<< m2 >>
rect 236 2980 280 3024
<< m3 >>
rect 236 2980 280 3024
<< via2 >>
rect 243 2987 273 3017
<< m2 >>
rect 819 1787 962 1817
<< m3 >>
rect 819 1787 849 2217
<< m2 >>
rect 819 2187 977 2217
<< m3 >>
rect 947 2187 977 2217
<< m2 >>
rect 371 2187 977 2217
<< m3 >>
rect 371 2187 401 2217
<< m2 >>
rect 243 2187 401 2217
<< m3 >>
rect 243 1787 273 2217
<< m2 >>
rect 243 1787 386 1817
<< m1 >>
rect 365 1777 411 1831
<< m2 >>
rect 365 1777 411 1831
<< via1 >>
rect 372 1784 404 1824
<< m1 >>
rect 941 1777 987 1831
<< m2 >>
rect 941 1777 987 1831
<< via1 >>
rect 948 1784 980 1824
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m2 >>
rect 812 1780 856 1824
<< m3 >>
rect 812 1780 856 1824
<< via2 >>
rect 819 1787 849 1817
<< m2 >>
rect 812 2180 856 2224
<< m3 >>
rect 812 2180 856 2224
<< via2 >>
rect 819 2187 849 2217
<< m2 >>
rect 940 2180 984 2224
<< m3 >>
rect 940 2180 984 2224
<< via2 >>
rect 947 2187 977 2217
<< m2 >>
rect 940 2180 984 2224
<< m3 >>
rect 940 2180 984 2224
<< via2 >>
rect 947 2187 977 2217
<< m2 >>
rect 364 2180 408 2224
<< m3 >>
rect 364 2180 408 2224
<< via2 >>
rect 371 2187 401 2217
<< m2 >>
rect 364 2180 408 2224
<< m3 >>
rect 364 2180 408 2224
<< via2 >>
rect 371 2187 401 2217
<< m2 >>
rect 236 2180 280 2224
<< m3 >>
rect 236 2180 280 2224
<< via2 >>
rect 243 2187 273 2217
<< m2 >>
rect 236 1780 280 1824
<< m3 >>
rect 236 1780 280 1824
<< via2 >>
rect 243 1787 273 1817
<< m3 >>
rect 659 538 689 1657
<< m3 >>
rect 659 1627 689 1657
<< m3 >>
rect 659 1627 689 2057
<< m3 >>
rect 659 2027 689 2057
<< m2 >>
rect 659 2027 1265 2057
<< m3 >>
rect 1235 2027 1265 2057
<< m3 >>
rect 1235 1642 1265 2057
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 1197 1617 1307 1671
<< m2 >>
rect 1197 1617 1307 1671
<< via1 >>
rect 1204 1624 1300 1664
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 621 517 731 571
<< m2 >>
rect 621 517 731 571
<< via1 >>
rect 628 524 724 564
<< m2 >>
rect 652 2020 696 2064
<< m3 >>
rect 652 2020 696 2064
<< via2 >>
rect 659 2027 689 2057
<< m2 >>
rect 1228 2020 1272 2064
<< m3 >>
rect 1228 2020 1272 2064
<< via2 >>
rect 1235 2027 1265 2057
<< m2 >>
rect 387 685 978 715
<< m3 >>
rect 948 685 978 715
<< m3 >>
rect 948 525 978 715
<< m2 >>
rect 948 525 1266 555
<< m3 >>
rect 1236 525 1266 555
<< m2 >>
rect 1236 525 1410 555
<< m3 >>
rect 1380 525 1410 2459
<< m2 >>
rect 1236 2429 1410 2459
<< m3 >>
rect 1236 2429 1266 2459
<< m3 >>
rect 1236 2429 1266 2859
<< m3 >>
rect 1236 2829 1266 2859
<< m2 >>
rect 660 2829 1266 2859
<< m3 >>
rect 660 2829 690 2859
<< m3 >>
rect 660 2444 690 2859
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 621 2417 731 2471
<< m2 >>
rect 621 2417 731 2471
<< via1 >>
rect 628 2424 724 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m2 >>
rect 941 678 985 722
<< m3 >>
rect 941 678 985 722
<< via2 >>
rect 948 685 978 715
<< m2 >>
rect 941 518 985 562
<< m3 >>
rect 941 518 985 562
<< via2 >>
rect 948 525 978 555
<< m2 >>
rect 1229 518 1273 562
<< m3 >>
rect 1229 518 1273 562
<< via2 >>
rect 1236 525 1266 555
<< m2 >>
rect 1229 518 1273 562
<< m3 >>
rect 1229 518 1273 562
<< via2 >>
rect 1236 525 1266 555
<< m2 >>
rect 1373 518 1417 562
<< m3 >>
rect 1373 518 1417 562
<< via2 >>
rect 1380 525 1410 555
<< m2 >>
rect 1373 2422 1417 2466
<< m3 >>
rect 1373 2422 1417 2466
<< via2 >>
rect 1380 2429 1410 2459
<< m2 >>
rect 1229 2422 1273 2466
<< m3 >>
rect 1229 2422 1273 2466
<< via2 >>
rect 1236 2429 1266 2459
<< m2 >>
rect 1229 2822 1273 2866
<< m3 >>
rect 1229 2822 1273 2866
<< via2 >>
rect 1236 2829 1266 2859
<< m2 >>
rect 653 2822 697 2866
<< m3 >>
rect 653 2822 697 2866
<< via2 >>
rect 660 2829 690 2859
<< m2 >>
rect 1251 3221 1410 3251
<< m3 >>
rect 1380 2709 1410 3251
<< m2 >>
rect 1044 2709 1410 2739
<< m3 >>
rect 1044 2709 1074 2739
<< m2 >>
rect 1044 2709 1506 2739
<< m3 >>
rect 1476 2309 1506 2739
<< m2 >>
rect 1044 2309 1506 2339
<< m3 >>
rect 1044 2309 1074 2339
<< m2 >>
rect 1044 2309 1506 2339
<< m3 >>
rect 1476 1909 1506 2339
<< m2 >>
rect 1044 1909 1506 1939
<< m3 >>
rect 1044 1909 1074 1939
<< m2 >>
rect 468 1909 1074 1939
<< m3 >>
rect 468 1909 498 1939
<< m2 >>
rect 148 1909 498 1939
<< m3 >>
rect 148 1909 178 2339
<< m2 >>
rect 148 2309 498 2339
<< m3 >>
rect 468 2309 498 2339
<< m2 >>
rect 148 2309 498 2339
<< m3 >>
rect 148 2309 178 2739
<< m2 >>
rect 148 2709 498 2739
<< m3 >>
rect 468 2709 498 2739
<< m2 >>
rect 148 2709 498 2739
<< m3 >>
rect 148 2709 178 3139
<< m2 >>
rect 148 3109 498 3139
<< m3 >>
rect 468 3109 498 3139
<< m2 >>
rect 468 3109 1059 3139
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 1005 3097 1115 3151
<< m2 >>
rect 1005 3097 1115 3151
<< via1 >>
rect 1012 3104 1108 3144
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 1197 3217 1307 3271
<< m2 >>
rect 1197 3217 1307 3271
<< via1 >>
rect 1204 3224 1300 3264
<< m2 >>
rect 1373 3214 1417 3258
<< m3 >>
rect 1373 3214 1417 3258
<< via2 >>
rect 1380 3221 1410 3251
<< m2 >>
rect 1373 2702 1417 2746
<< m3 >>
rect 1373 2702 1417 2746
<< via2 >>
rect 1380 2709 1410 2739
<< m2 >>
rect 1037 2702 1081 2746
<< m3 >>
rect 1037 2702 1081 2746
<< via2 >>
rect 1044 2709 1074 2739
<< m2 >>
rect 1037 2702 1081 2746
<< m3 >>
rect 1037 2702 1081 2746
<< via2 >>
rect 1044 2709 1074 2739
<< m2 >>
rect 1469 2702 1513 2746
<< m3 >>
rect 1469 2702 1513 2746
<< via2 >>
rect 1476 2709 1506 2739
<< m2 >>
rect 1469 2302 1513 2346
<< m3 >>
rect 1469 2302 1513 2346
<< via2 >>
rect 1476 2309 1506 2339
<< m2 >>
rect 1037 2302 1081 2346
<< m3 >>
rect 1037 2302 1081 2346
<< via2 >>
rect 1044 2309 1074 2339
<< m2 >>
rect 1037 2302 1081 2346
<< m3 >>
rect 1037 2302 1081 2346
<< via2 >>
rect 1044 2309 1074 2339
<< m2 >>
rect 1469 2302 1513 2346
<< m3 >>
rect 1469 2302 1513 2346
<< via2 >>
rect 1476 2309 1506 2339
<< m2 >>
rect 1469 1902 1513 1946
<< m3 >>
rect 1469 1902 1513 1946
<< via2 >>
rect 1476 1909 1506 1939
<< m2 >>
rect 1037 1902 1081 1946
<< m3 >>
rect 1037 1902 1081 1946
<< via2 >>
rect 1044 1909 1074 1939
<< m2 >>
rect 1037 1902 1081 1946
<< m3 >>
rect 1037 1902 1081 1946
<< via2 >>
rect 1044 1909 1074 1939
<< m2 >>
rect 461 1902 505 1946
<< m3 >>
rect 461 1902 505 1946
<< via2 >>
rect 468 1909 498 1939
<< m2 >>
rect 461 1902 505 1946
<< m3 >>
rect 461 1902 505 1946
<< via2 >>
rect 468 1909 498 1939
<< m2 >>
rect 141 1902 185 1946
<< m3 >>
rect 141 1902 185 1946
<< via2 >>
rect 148 1909 178 1939
<< m2 >>
rect 141 2302 185 2346
<< m3 >>
rect 141 2302 185 2346
<< via2 >>
rect 148 2309 178 2339
<< m2 >>
rect 461 2302 505 2346
<< m3 >>
rect 461 2302 505 2346
<< via2 >>
rect 468 2309 498 2339
<< m2 >>
rect 461 2302 505 2346
<< m3 >>
rect 461 2302 505 2346
<< via2 >>
rect 468 2309 498 2339
<< m2 >>
rect 141 2302 185 2346
<< m3 >>
rect 141 2302 185 2346
<< via2 >>
rect 148 2309 178 2339
<< m2 >>
rect 141 2702 185 2746
<< m3 >>
rect 141 2702 185 2746
<< via2 >>
rect 148 2709 178 2739
<< m2 >>
rect 461 2702 505 2746
<< m3 >>
rect 461 2702 505 2746
<< via2 >>
rect 468 2709 498 2739
<< m2 >>
rect 461 2702 505 2746
<< m3 >>
rect 461 2702 505 2746
<< via2 >>
rect 468 2709 498 2739
<< m2 >>
rect 141 2702 185 2746
<< m3 >>
rect 141 2702 185 2746
<< via2 >>
rect 148 2709 178 2739
<< m2 >>
rect 141 3102 185 3146
<< m3 >>
rect 141 3102 185 3146
<< via2 >>
rect 148 3109 178 3139
<< m2 >>
rect 461 3102 505 3146
<< m3 >>
rect 461 3102 505 3146
<< via2 >>
rect 468 3109 498 3139
<< m2 >>
rect 461 3102 505 3146
<< m3 >>
rect 461 3102 505 3146
<< via2 >>
rect 468 3109 498 3139
<< m2 >>
rect 1154 9002 2177 9032
<< m3 >>
rect 1154 3386 1184 9032
<< m2 >>
rect 946 3386 1184 3416
<< m3 >>
rect 946 3386 976 3416
<< m3 >>
rect 946 3226 976 3416
<< m2 >>
rect 673 3226 976 3256
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 621 3217 731 3271
<< m2 >>
rect 621 3217 731 3271
<< via1 >>
rect 628 3224 724 3264
<< locali >>
rect 2103 8957 2261 9091
<< m1 >>
rect 2103 8957 2261 9091
<< viali >>
rect 2110 8964 2254 9084
<< m2 >>
rect 1147 8995 1191 9039
<< m3 >>
rect 1147 8995 1191 9039
<< via2 >>
rect 1154 9002 1184 9032
<< m2 >>
rect 1147 3379 1191 3423
<< m3 >>
rect 1147 3379 1191 3423
<< via2 >>
rect 1154 3386 1184 3416
<< m2 >>
rect 939 3379 983 3423
<< m3 >>
rect 939 3379 983 3423
<< via2 >>
rect 946 3386 976 3416
<< m2 >>
rect 939 3219 983 3263
<< m3 >>
rect 939 3219 983 3263
<< via2 >>
rect 946 3226 976 3256
<< m3 >>
rect 434 7499 464 9018
<< m2 >>
rect 434 7499 2192 7529
<< m3 >>
rect 2162 7242 2192 7529
<< locali >>
rect 375 8957 533 9091
<< m1 >>
rect 375 8957 533 9091
<< viali >>
rect 382 8964 526 9084
<< locali >>
rect 2103 7177 2261 7311
<< m1 >>
rect 2103 7177 2261 7311
<< viali >>
rect 2110 7184 2254 7304
<< m2 >>
rect 427 7492 471 7536
<< m3 >>
rect 427 7492 471 7536
<< via2 >>
rect 434 7499 464 7529
<< m2 >>
rect 2155 7492 2199 7536
<< m3 >>
rect 2155 7492 2199 7536
<< via2 >>
rect 2162 7499 2192 7529
<< m3 >>
rect 434 6249 464 7240
<< m2 >>
rect 434 6249 2192 6279
<< m3 >>
rect 2162 5464 2192 6279
<< locali >>
rect 375 7177 533 7311
<< m1 >>
rect 375 7177 533 7311
<< viali >>
rect 382 7184 526 7304
<< locali >>
rect 2103 5407 2261 5541
<< m1 >>
rect 2103 5407 2261 5541
<< viali >>
rect 2110 5414 2254 5534
<< m2 >>
rect 427 6242 471 6286
<< m3 >>
rect 427 6242 471 6286
<< via2 >>
rect 434 6249 464 6279
<< m2 >>
rect 2155 6242 2199 6286
<< m3 >>
rect 2155 6242 2199 6286
<< via2 >>
rect 2162 6249 2192 6279
<< locali >>
rect 100 9274 2536 9324
<< locali >>
rect 100 100 2536 150
<< m1 >>
rect 100 150 150 9274
<< m1 >>
rect 2486 150 2536 9274
<< locali >>
rect 93 9267 157 9331
<< m1 >>
rect 93 9267 157 9331
<< viali >>
rect 100 9274 150 9324
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2479 9267 2543 9331
<< m1 >>
rect 2479 9267 2543 9331
<< viali >>
rect 2486 9274 2536 9324
<< locali >>
rect 2479 93 2543 157
<< m1 >>
rect 2479 93 2543 157
<< viali >>
rect 2486 100 2536 150
<< locali >>
rect 0 9374 2636 9424
<< locali >>
rect 0 0 2636 50
<< m1 >>
rect 0 50 50 9374
<< m1 >>
rect 2586 50 2636 9374
<< locali >>
rect -7 9367 57 9431
<< m1 >>
rect -7 9367 57 9431
<< viali >>
rect 0 9374 50 9424
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2579 9367 2643 9431
<< m1 >>
rect 2579 9367 2643 9431
<< viali >>
rect 2586 9374 2636 9424
<< locali >>
rect 2579 -7 2643 57
<< m1 >>
rect 2579 -7 2643 57
<< viali >>
rect 2586 0 2636 50
<< locali >>
rect 208 5414 526 5534
<< locali >>
rect 100 9168 2536 9224
<< locali >>
rect 93 9161 157 9231
<< m1 >>
rect 93 9161 157 9231
<< viali >>
rect 100 9168 150 9224
<< locali >>
rect 2479 9161 2543 9231
<< m1 >>
rect 2479 9161 2543 9231
<< viali >>
rect 2486 9168 2536 9224
<< locali >>
rect 100 7504 2536 7560
<< locali >>
rect 93 7497 157 7567
<< m1 >>
rect 93 7497 157 7567
<< viali >>
rect 100 7504 150 7560
<< locali >>
rect 2479 7497 2543 7567
<< m1 >>
rect 2479 7497 2543 7567
<< viali >>
rect 2486 7504 2536 7560
<< locali >>
rect 100 7388 2536 7444
<< locali >>
rect 93 7381 157 7451
<< m1 >>
rect 93 7381 157 7451
<< viali >>
rect 100 7388 150 7444
<< locali >>
rect 2479 7381 2543 7451
<< m1 >>
rect 2479 7381 2543 7451
<< viali >>
rect 2486 7388 2536 7444
<< locali >>
rect 100 5724 2536 5780
<< locali >>
rect 93 5717 157 5787
<< m1 >>
rect 93 5717 157 5787
<< viali >>
rect 100 5724 150 5780
<< locali >>
rect 2479 5717 2543 5787
<< m1 >>
rect 2479 5717 2543 5787
<< viali >>
rect 2486 5724 2536 5780
<< locali >>
rect 100 5618 2536 5674
<< locali >>
rect 93 5611 157 5681
<< m1 >>
rect 93 5611 157 5681
<< viali >>
rect 100 5618 150 5674
<< locali >>
rect 2479 5611 2543 5681
<< m1 >>
rect 2479 5611 2543 5681
<< viali >>
rect 2486 5618 2536 5674
<< locali >>
rect 100 3954 2536 4010
<< locali >>
rect 93 3947 157 4017
<< m1 >>
rect 93 3947 157 4017
<< viali >>
rect 100 3954 150 4010
<< locali >>
rect 2479 3947 2543 4017
<< m1 >>
rect 2479 3947 2543 4017
<< viali >>
rect 2486 3954 2536 4010
<< locali >>
rect 820 3504 1108 3544
<< locali >>
rect 244 3504 532 3544
<< locali >>
rect 628 3384 788 3424
<< locali >>
rect 820 804 1108 844
<< locali >>
rect 1204 684 1364 724
<< locali >>
rect 244 804 532 844
<< locali >>
rect 0 1436 2636 1532
<< locali >>
rect -7 1429 57 1539
<< m1 >>
rect -7 1429 57 1539
<< viali >>
rect 0 1436 50 1532
<< locali >>
rect 2579 1429 2643 1539
<< m1 >>
rect 2579 1429 2643 1539
<< viali >>
rect 2586 1436 2636 1532
<< locali >>
rect 0 3676 2636 3772
<< locali >>
rect -7 3669 57 3779
<< m1 >>
rect -7 3669 57 3779
<< viali >>
rect 0 3676 50 3772
<< locali >>
rect 2579 3669 2643 3779
<< m1 >>
rect 2579 3669 2643 3779
<< viali >>
rect 2586 3676 2636 3772
<< locali >>
rect 100 976 2536 1072
<< locali >>
rect 93 969 157 1079
<< m1 >>
rect 93 969 157 1079
<< viali >>
rect 100 976 150 1072
<< locali >>
rect 2479 969 2543 1079
<< m1 >>
rect 2479 969 2543 1079
<< viali >>
rect 2486 976 2536 1072
<< locali >>
rect 100 336 2536 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< locali >>
rect 2479 329 2543 439
<< m1 >>
rect 2479 329 2543 439
<< viali >>
rect 2486 336 2536 432
<< labels >>
flabel m2 s 819 2987 962 3017 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 819 1787 962 1817 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 0 9374 2636 9424 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 100 9274 2536 9324 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m3 s 659 538 689 1657 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744372385
<< checkpaint >>
rect 0 0 0 0
<< labels >>
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1746459945
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 14358 5948 14408
<< locali >>
rect -100 -100 5948 -50
<< m1 >>
rect -100 -50 -50 14358
<< m1 >>
rect 5898 -50 5948 14358
<< locali >>
rect -107 14351 -43 14415
<< m1 >>
rect -107 14351 -43 14415
<< viali >>
rect -100 14358 -50 14408
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 5891 14351 5955 14415
<< m1 >>
rect 5891 14351 5955 14415
<< viali >>
rect 5898 14358 5948 14408
<< locali >>
rect 5891 -107 5955 -43
<< m1 >>
rect 5891 -107 5955 -43
<< viali >>
rect 5898 -100 5948 -50
<< locali >>
rect -200 14458 6048 14508
<< locali >>
rect -200 -200 6048 -150
<< m1 >>
rect -200 -150 -150 14458
<< m1 >>
rect 5998 -150 6048 14458
<< locali >>
rect -207 14451 -143 14515
<< m1 >>
rect -207 14451 -143 14515
<< viali >>
rect -200 14458 -150 14508
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 5991 14451 6055 14515
<< m1 >>
rect 5991 14451 6055 14515
<< viali >>
rect 5998 14458 6048 14508
<< locali >>
rect 5991 -207 6055 -143
<< m1 >>
rect 5991 -207 6055 -143
<< viali >>
rect 5998 -200 6048 -150
use JNW_GR06 U1_JNW_GR06 
transform 1 0 0 0 1 0
box 0 0 1390 8118
<< labels >>
flabel locali s -200 14458 6048 14508 0 FreeSans 400 0 0 0 VDD
port 205 nsew signal bidirectional
flabel locali s -100 14358 5948 14408 0 FreeSans 400 0 0 0 VSS
port 206 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1745941688
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 500
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 260
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 500
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 260
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 900
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP3<1>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 1300
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 900
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP3<0>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 1300
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 3700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 3700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 3300
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4<1>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 3060
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 3300
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4<0>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 3060
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 4100
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 4500
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 4100
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 4500
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 2100
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 2500
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 3512 0 1 1860
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 2100
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 2500
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2936 0 1 1860
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2320
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4170
box 0 0 2236 1720
use AALMISC_CAP50f None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 4488 0 1 500
box 0 0 580 842
<< locali >>
rect 100 6240 5268 6290
<< locali >>
rect 100 100 5268 150
<< m1 >>
rect 100 150 150 6240
<< m1 >>
rect 5218 150 5268 6240
<< locali >>
rect 93 6233 157 6297
<< m1 >>
rect 93 6233 157 6297
<< viali >>
rect 100 6240 150 6290
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 5211 6233 5275 6297
<< m1 >>
rect 5211 6233 5275 6297
<< viali >>
rect 5218 6240 5268 6290
<< locali >>
rect 5211 93 5275 157
<< m1 >>
rect 5211 93 5275 157
<< viali >>
rect 5218 100 5268 150
<< locali >>
rect 0 6340 5368 6390
<< locali >>
rect 0 0 5368 50
<< m1 >>
rect 0 50 50 6340
<< m1 >>
rect 5318 50 5368 6340
<< locali >>
rect -7 6333 57 6397
<< m1 >>
rect -7 6333 57 6397
<< viali >>
rect 0 6340 50 6390
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 5311 6333 5375 6397
<< m1 >>
rect 5311 6333 5375 6397
<< viali >>
rect 5318 6340 5368 6390
<< locali >>
rect 5311 -7 5375 57
<< m1 >>
rect 5311 -7 5375 57
<< viali >>
rect 5318 0 5368 50
<< locali >>
rect 2888 4400 3176 4440
<< locali >>
rect 3464 4400 3752 4440
<< locali >>
rect 3848 4280 4008 4320
<< locali >>
rect 3464 2400 3752 2440
<< locali >>
rect 3848 2280 4008 2320
<< locali >>
rect 2888 2400 3176 2440
<< locali >>
rect 2736 332 3712 428
<< locali >>
rect 2729 325 2793 435
<< m1 >>
rect 2729 325 2793 435
<< viali >>
rect 2736 332 2786 428
<< locali >>
rect 3655 325 3719 435
<< m1 >>
rect 3655 325 3719 435
<< viali >>
rect 3662 332 3712 428
<< locali >>
rect 3312 1372 4288 1468
<< locali >>
rect 3305 1365 3369 1475
<< m1 >>
rect 3305 1365 3369 1475
<< viali >>
rect 3312 1372 3362 1468
<< locali >>
rect 4231 1365 4295 1475
<< m1 >>
rect 4231 1365 4295 1475
<< viali >>
rect 4238 1372 4288 1468
<< locali >>
rect 2736 3132 3712 3228
<< locali >>
rect 2729 3125 2793 3235
<< m1 >>
rect 2729 3125 2793 3235
<< viali >>
rect 2736 3132 2786 3228
<< locali >>
rect 3655 3125 3719 3235
<< m1 >>
rect 3655 3125 3719 3235
<< viali >>
rect 3662 3132 3712 3228
<< locali >>
rect 2736 4572 3712 4668
<< locali >>
rect 2729 4565 2793 4675
<< m1 >>
rect 2729 4565 2793 4675
<< viali >>
rect 2736 4572 2786 4668
<< locali >>
rect 3655 4565 3719 4675
<< m1 >>
rect 3655 4565 3719 4675
<< viali >>
rect 3662 4572 3712 4668
<< locali >>
rect 3312 2572 4288 2668
<< locali >>
rect 3305 2565 3369 2675
<< m1 >>
rect 3305 2565 3369 2675
<< viali >>
rect 3312 2572 3362 2668
<< locali >>
rect 4231 2565 4295 2675
<< m1 >>
rect 4231 2565 4295 2675
<< viali >>
rect 4238 2572 4288 2668
<< locali >>
rect 3312 1932 4288 2028
<< locali >>
rect 3305 1925 3369 2035
<< m1 >>
rect 3305 1925 3369 2035
<< viali >>
rect 3312 1932 3362 2028
<< locali >>
rect 4231 1925 4295 2035
<< m1 >>
rect 4231 1925 4295 2035
<< viali >>
rect 4238 1932 4288 2028
<< locali >>
rect 308 5630 626 5750
<< locali >>
rect 0 2164 5368 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 5311 2157 5375 2227
<< m1 >>
rect 5311 2157 5375 2227
<< viali >>
rect 5318 2164 5368 2220
<< locali >>
rect 0 500 5368 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 5311 493 5375 563
<< m1 >>
rect 5311 493 5375 563
<< viali >>
rect 5318 500 5368 556
<< locali >>
rect 0 3984 5368 4040
<< locali >>
rect -7 3977 57 4047
<< m1 >>
rect -7 3977 57 4047
<< viali >>
rect 0 3984 50 4040
<< locali >>
rect 5311 3977 5375 4047
<< m1 >>
rect 5311 3977 5375 4047
<< viali >>
rect 5318 3984 5368 4040
<< locali >>
rect 0 2320 5368 2376
<< locali >>
rect -7 2313 57 2383
<< m1 >>
rect -7 2313 57 2383
<< viali >>
rect 0 2320 50 2376
<< locali >>
rect 5311 2313 5375 2383
<< m1 >>
rect 5311 2313 5375 2383
<< viali >>
rect 5318 2320 5368 2376
<< locali >>
rect 0 5834 5368 5890
<< locali >>
rect -7 5827 57 5897
<< m1 >>
rect -7 5827 57 5897
<< viali >>
rect 0 5834 50 5890
<< locali >>
rect 5311 5827 5375 5897
<< m1 >>
rect 5311 5827 5375 5897
<< viali >>
rect 5318 5834 5368 5890
<< locali >>
rect 0 4170 5368 4226
<< locali >>
rect -7 4163 57 4233
<< m1 >>
rect -7 4163 57 4233
<< viali >>
rect 0 4170 50 4226
<< locali >>
rect 5311 4163 5375 4233
<< m1 >>
rect 5311 4163 5375 4233
<< viali >>
rect 5318 4170 5368 4226
<< labels >>
flabel locali s 100 6240 5268 6290 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 0 6340 5368 6390 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
<< properties >>
<< end >>
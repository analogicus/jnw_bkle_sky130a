magic
tech sky130A
magscale 1 1
timestamp 1726667330
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 x1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 0 0
rect 0 0 0 0
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 0 0
<< labels >>
<< properties >>
<< end >>
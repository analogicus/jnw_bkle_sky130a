magic
tech sky130A
magscale 1 1
timestamp 1745323676
<< checkpaint >>
rect 0 0 1000 1000
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6460
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWTR_CAPX1 None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 540 540
use JNWATR_PCH_4C5F0 None_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7800 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7224 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7800 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7224 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7800 0 1 6700
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7224 0 1 7000
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7800 0 1 7000
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN1<2>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7800 0 1 7400
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN1<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6700
box 0 0 576 400
use JNWTR_RPPO8 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 1820
box 0 0 1372 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4280
box 0 0 940 1720
use AALMISC_PNP_W3p40L3p40 load1_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 8080
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<0> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<1> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<2> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<3> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<4> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<5> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<6> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
use AALMISC_PNP_W3p40L3p40 load1_QP2<7> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6700
box 0 0 1340 1340
<< locali >>
rect 100 9770 8576 9820
<< locali >>
rect 100 100 8576 150
<< m1 >>
rect 100 150 150 9770
<< m1 >>
rect 8526 150 8576 9770
<< locali >>
rect 93 9763 157 9827
<< m1 >>
rect 93 9763 157 9827
<< viali >>
rect 100 9770 150 9820
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 8519 9763 8583 9827
<< m1 >>
rect 8519 9763 8583 9827
<< viali >>
rect 8526 9770 8576 9820
<< locali >>
rect 8519 93 8583 157
<< m1 >>
rect 8519 93 8583 157
<< viali >>
rect 8526 100 8576 150
<< locali >>
rect 0 9870 8676 9920
<< locali >>
rect 0 0 8676 50
<< m1 >>
rect 0 50 50 9870
<< m1 >>
rect 8626 50 8676 9870
<< locali >>
rect -7 9863 57 9927
<< m1 >>
rect -7 9863 57 9927
<< viali >>
rect 0 9870 50 9920
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 8619 9863 8683 9927
<< m1 >>
rect 8619 9863 8683 9927
<< viali >>
rect 8626 9870 8676 9920
<< locali >>
rect 8619 -7 8683 57
<< m1 >>
rect 8619 -7 8683 57
<< viali >>
rect 8626 0 8676 50
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 7752 7000 8040 7040
<< locali >>
rect 8136 6880 8296 6920
<< locali >>
rect 7176 7000 7464 7040
<< locali >>
rect 7560 6880 7720 6920
<< locali >>
rect 7752 7000 8040 7040
<< locali >>
rect 8136 6880 8296 6920
<< locali >>
rect 7176 7000 7464 7040
<< locali >>
rect 7560 6880 7720 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 7752 7000 8040 7040
<< locali >>
rect 8136 6880 8296 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 7176 7300 7464 7340
<< locali >>
rect 7560 7180 7720 7220
<< locali >>
rect 7752 7300 8040 7340
<< locali >>
rect 8136 7180 8296 7220
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 636 6880 796 6920
<< locali >>
rect 252 7000 540 7040
<< locali >>
rect 100 6532 8576 6628
<< locali >>
rect 93 6525 157 6635
<< m1 >>
rect 93 6525 157 6635
<< viali >>
rect 100 6532 150 6628
<< locali >>
rect 8519 6525 8583 6635
<< m1 >>
rect 8519 6525 8583 6635
<< viali >>
rect 8526 6532 8576 6628
use OTA U1_OTA 
transform 1 0 2886 0 1 0
box 0 0 2886 11510
<< labels >>
flabel locali s 100 9770 8576 9820 0 FreeSans 400 0 0 0 VDD
port 36 nsew signal bidirectional
flabel locali s 0 9870 8676 9920 0 FreeSans 400 0 0 0 VSS
port 37 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744112857
<< checkpaint >>
rect 0 0 0 0
use JNWATR_PCH_4C1F2 diff1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 1600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT diff1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 1360
box 0 0 576 240
use JNWATR_PCH_4C1F2 diff1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 1600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT diff1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 1360
box 0 0 576 240
use JNWATR_PCH_4C5F0 mirror1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 2000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP mirror1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 2400
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror3_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 0
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror3_MN4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 -240
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror4_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror4_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 800
box 0 0 576 240
use JNWATR_PCH_4C5F0 mirror1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP mirror1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2400
box 0 0 576 240
use JNWATR_PCH_12C5F0 mirror1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 3200
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP mirror1_MP3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 3600
box 0 0 832 240
use JNWATR_PCH_12CTAPBOT mirror1_MP3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2960
box 0 0 832 240
use JNWATR_NCH_4C5F0 mirror4_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror4_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 800
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror3_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 0
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror3_MN3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 -240
box 0 0 576 240
use JNWATR_PCH_12C5F0 mirror1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 3200
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP mirror1_MP4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 3600
box 0 0 832 240
use JNWATR_PCH_12CTAPBOT mirror1_MP4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 2960
box 0 0 832 240
use JNWTR_RPPO2 None_R1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 2496 0 1 400
box 0 0 724 1720
use JNWTR_RPPO2 None_R2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 0 0 1 400
box 0 0 724 1720
<< locali >>
rect -250 3950 3470 4050
<< locali >>
rect -250 -450 3470 -350
<< m1 >>
rect -250 -350 -150 3950
<< m1 >>
rect 3370 -350 3470 3950
<< locali >>
rect -257 3943 -143 4057
<< m1 >>
rect -257 3943 -143 4057
<< viali >>
rect -250 3950 -150 4050
<< locali >>
rect -257 -457 -143 -343
<< m1 >>
rect -257 -457 -143 -343
<< viali >>
rect -250 -450 -150 -350
<< locali >>
rect 3363 3943 3477 4057
<< m1 >>
rect 3363 3943 3477 4057
<< viali >>
rect 3370 3950 3470 4050
<< locali >>
rect 3363 -457 3477 -343
<< m1 >>
rect 3363 -457 3477 -343
<< viali >>
rect 3370 -450 3470 -350
<< locali >>
rect -400 4100 3620 4200
<< locali >>
rect -400 -600 3620 -500
<< m1 >>
rect -400 -500 -300 4100
<< m1 >>
rect 3520 -500 3620 4100
<< locali >>
rect -407 4093 -293 4207
<< m1 >>
rect -407 4093 -293 4207
<< viali >>
rect -400 4100 -300 4200
<< locali >>
rect -407 -607 -293 -493
<< m1 >>
rect -407 -607 -293 -493
<< viali >>
rect -400 -600 -300 -500
<< locali >>
rect 3513 4093 3627 4207
<< m1 >>
rect 3513 4093 3627 4207
<< viali >>
rect 3520 4100 3620 4200
<< locali >>
rect 3513 -607 3627 -493
<< m1 >>
rect 3513 -607 3627 -493
<< viali >>
rect 3520 -600 3620 -500
<< locali >>
rect 1040 2300 1328 2340
<< locali >>
rect 1040 300 1328 340
<< locali >>
rect 1040 700 1328 740
<< locali >>
rect 1616 2300 1904 2340
<< locali >>
rect 2000 2180 2160 2220
<< locali >>
rect 1616 3500 1904 3540
<< locali >>
rect 2256 3380 2416 3420
<< locali >>
rect 1616 700 1904 740
<< locali >>
rect 2000 580 2160 620
<< locali >>
rect 1616 300 1904 340
<< locali >>
rect 2000 180 2160 220
<< locali >>
rect 784 3500 1072 3540
<< locali >>
rect -250 1432 3470 1528
<< locali >>
rect -257 1425 -143 1535
<< m1 >>
rect -257 1425 -143 1535
<< viali >>
rect -250 1432 -150 1528
<< locali >>
rect 3363 1425 3477 1535
<< m1 >>
rect 3363 1425 3477 1535
<< viali >>
rect 3370 1432 3470 1528
<< locali >>
rect -250 2472 3470 2568
<< locali >>
rect -257 2465 -143 2575
<< m1 >>
rect -257 2465 -143 2575
<< viali >>
rect -250 2472 -150 2568
<< locali >>
rect 3363 2465 3477 2575
<< m1 >>
rect 3363 2465 3477 2575
<< viali >>
rect 3370 2472 3470 2568
<< locali >>
rect -400 -168 3620 -72
<< locali >>
rect -407 -175 -293 -65
<< m1 >>
rect -407 -175 -293 -65
<< viali >>
rect -400 -168 -300 -72
<< locali >>
rect 3513 -175 3627 -65
<< m1 >>
rect 3513 -175 3627 -65
<< viali >>
rect 3520 -168 3620 -72
<< locali >>
rect -400 872 3620 968
<< locali >>
rect -407 865 -293 975
<< m1 >>
rect -407 865 -293 975
<< viali >>
rect -400 872 -300 968
<< locali >>
rect 3513 865 3627 975
<< m1 >>
rect 3513 865 3627 975
<< viali >>
rect 3520 872 3620 968
<< locali >>
rect -250 3672 3470 3768
<< locali >>
rect -257 3665 -143 3775
<< m1 >>
rect -257 3665 -143 3775
<< viali >>
rect -250 3672 -150 3768
<< locali >>
rect 3363 3665 3477 3775
<< m1 >>
rect 3363 3665 3477 3775
<< viali >>
rect 3370 3672 3470 3768
<< locali >>
rect -250 3032 3470 3128
<< locali >>
rect -257 3025 -143 3135
<< m1 >>
rect -257 3025 -143 3135
<< viali >>
rect -250 3032 -150 3128
<< locali >>
rect 3363 3025 3477 3135
<< m1 >>
rect 3363 3025 3477 3135
<< viali >>
rect 3370 3032 3470 3128
<< labels >>
flabel locali s -250 3950 3470 4050 0 FreeSans 400 0 0 0 VDD
port 8 nsew signal bidirectional
flabel locali s -400 4100 3620 4200 0 FreeSans 400 0 0 0 VSS
port 9 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1745089113
<< checkpaint >>
rect 0 0 0 0
<< locali >>
rect -100 9090 8070 9140
<< locali >>
rect -100 -100 8070 -50
<< m1 >>
rect -100 -50 -50 9090
<< m1 >>
rect 8020 -50 8070 9090
<< locali >>
rect -107 9083 -43 9147
<< m1 >>
rect -107 9083 -43 9147
<< viali >>
rect -100 9090 -50 9140
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 8013 9083 8077 9147
<< m1 >>
rect 8013 9083 8077 9147
<< viali >>
rect 8020 9090 8070 9140
<< locali >>
rect 8013 -107 8077 -43
<< m1 >>
rect 8013 -107 8077 -43
<< viali >>
rect 8020 -100 8070 -50
<< locali >>
rect -200 9190 8170 9240
<< locali >>
rect -200 -200 8170 -150
<< m1 >>
rect -200 -150 -150 9190
<< m1 >>
rect 8120 -150 8170 9190
<< locali >>
rect -207 9183 -143 9247
<< m1 >>
rect -207 9183 -143 9247
<< viali >>
rect -200 9190 -150 9240
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 8113 9183 8177 9247
<< m1 >>
rect 8113 9183 8177 9247
<< viali >>
rect 8120 9190 8170 9240
<< locali >>
rect 8113 -207 8177 -143
<< m1 >>
rect 8113 -207 8177 -143
<< viali >>
rect 8120 -200 8170 -150
use JNW_GR06 U1_JNW_GR06 
transform 1 0 0 0 1 0
box 0 0 2714 6290
<< labels >>
flabel locali s -100 9090 8070 9140 0 FreeSans 400 0 0 0 VDD
port 51 nsew signal bidirectional
flabel locali s -200 9190 8170 9240 0 FreeSans 400 0 0 0 VSS
port 52 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744380266
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1400
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1160
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1400
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 2760
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 2760
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3400
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 3400
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 600
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1000
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT mirror2_MN4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 360
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 600
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1000
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT mirror2_MN3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 360
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 2200
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 1800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 2200
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 3800
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 4200
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 3800
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2128 0 1 4200
box 0 0 576 240
<< locali >>
rect 150 4550 2954 4650
<< locali >>
rect 150 150 2954 250
<< m1 >>
rect 150 250 250 4550
<< m1 >>
rect 2854 250 2954 4550
<< locali >>
rect 143 4543 257 4657
<< m1 >>
rect 143 4543 257 4657
<< viali >>
rect 150 4550 250 4650
<< locali >>
rect 143 143 257 257
<< m1 >>
rect 143 143 257 257
<< viali >>
rect 150 150 250 250
<< locali >>
rect 2847 4543 2961 4657
<< m1 >>
rect 2847 4543 2961 4657
<< viali >>
rect 2854 4550 2954 4650
<< locali >>
rect 2847 143 2961 257
<< m1 >>
rect 2847 143 2961 257
<< viali >>
rect 2854 150 2954 250
<< locali >>
rect 0 4700 3104 4800
<< locali >>
rect 0 0 3104 100
<< m1 >>
rect 0 100 100 4700
<< m1 >>
rect 3004 100 3104 4700
<< locali >>
rect -7 4693 107 4807
<< m1 >>
rect -7 4693 107 4807
<< viali >>
rect 0 4700 100 4800
<< locali >>
rect -7 -7 107 107
<< m1 >>
rect -7 -7 107 107
<< viali >>
rect 0 0 100 100
<< locali >>
rect 2997 4693 3111 4807
<< m1 >>
rect 2997 4693 3111 4807
<< viali >>
rect 3004 4700 3104 4800
<< locali >>
rect 2997 -7 3111 107
<< m1 >>
rect 2997 -7 3111 107
<< viali >>
rect 3004 0 3104 100
<< locali >>
rect 352 3300 640 3340
<< locali >>
rect 736 3180 896 3220
<< locali >>
rect 2080 3300 2368 3340
<< locali >>
rect 352 3700 640 3740
<< locali >>
rect 2080 3700 2368 3740
<< locali >>
rect 2464 3580 2624 3620
<< locali >>
rect 352 900 640 940
<< locali >>
rect 2080 900 2368 940
<< locali >>
rect 2464 780 2624 820
<< locali >>
rect 352 2100 640 2140
<< locali >>
rect 736 1980 896 2020
<< locali >>
rect 2080 2100 2368 2140
<< locali >>
rect 352 4100 640 4140
<< locali >>
rect 2080 4100 2368 4140
<< locali >>
rect 0 1232 3104 1328
<< locali >>
rect -7 1225 107 1335
<< m1 >>
rect -7 1225 107 1335
<< viali >>
rect 0 1232 100 1328
<< locali >>
rect 2997 1225 3111 1335
<< m1 >>
rect 2997 1225 3111 1335
<< viali >>
rect 3004 1232 3104 1328
<< locali >>
rect 150 2832 2954 2928
<< locali >>
rect 143 2825 257 2935
<< m1 >>
rect 143 2825 257 2935
<< viali >>
rect 150 2832 250 2928
<< locali >>
rect 2847 2825 2961 2935
<< m1 >>
rect 2847 2825 2961 2935
<< viali >>
rect 2854 2832 2954 2928
<< locali >>
rect 0 1072 3104 1168
<< locali >>
rect -7 1065 107 1175
<< m1 >>
rect -7 1065 107 1175
<< viali >>
rect 0 1072 100 1168
<< locali >>
rect 2997 1065 3111 1175
<< m1 >>
rect 2997 1065 3111 1175
<< viali >>
rect 3004 1072 3104 1168
<< locali >>
rect 0 432 3104 528
<< locali >>
rect -7 425 107 535
<< m1 >>
rect -7 425 107 535
<< viali >>
rect 0 432 100 528
<< locali >>
rect 2997 425 3111 535
<< m1 >>
rect 2997 425 3111 535
<< viali >>
rect 3004 432 3104 528
<< locali >>
rect 0 2272 3104 2368
<< locali >>
rect -7 2265 107 2375
<< m1 >>
rect -7 2265 107 2375
<< viali >>
rect 0 2272 100 2368
<< locali >>
rect 2997 2265 3111 2375
<< m1 >>
rect 2997 2265 3111 2375
<< viali >>
rect 3004 2272 3104 2368
<< locali >>
rect 150 4272 2954 4368
<< locali >>
rect 143 4265 257 4375
<< m1 >>
rect 143 4265 257 4375
<< viali >>
rect 150 4272 250 4368
<< locali >>
rect 2847 4265 2961 4375
<< m1 >>
rect 2847 4265 2961 4375
<< viali >>
rect 2854 4272 2954 4368
<< labels >>
flabel locali s 0 4700 3104 4800 0 FreeSans 400 0 0 0 VSS
port 43 nsew signal bidirectional
flabel locali s 150 4550 2954 4650 0 FreeSans 400 0 0 0 VDD
port 44 nsew signal bidirectional
<< properties >>
<< end >>
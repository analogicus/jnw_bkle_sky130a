magic
tech sky130A
magscale 1 1
timestamp 1745323676
<< checkpaint >>
rect 0 0 1000 1000
use JNWTR_RPPO4 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2920
box 0 0 940 1720
use JNWTR_RPPO4 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 5340
box 0 0 940 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 940 1720
use JNWTR_CAPX1 None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 7760
box 0 0 540 540
use JNWATR_NCH_2C1F2 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9000
box 0 0 512 400
use JNWATR_NCH_2CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9400
box 0 0 512 240
use JNWATR_NCH_2CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8760
box 0 0 512 240
<< locali >>
rect 100 9750 1440 9800
<< locali >>
rect 100 100 1440 150
<< m1 >>
rect 100 150 150 9750
<< m1 >>
rect 1390 150 1440 9750
<< locali >>
rect 93 9743 157 9807
<< m1 >>
rect 93 9743 157 9807
<< viali >>
rect 100 9750 150 9800
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1383 9743 1447 9807
<< m1 >>
rect 1383 9743 1447 9807
<< viali >>
rect 1390 9750 1440 9800
<< locali >>
rect 1383 93 1447 157
<< m1 >>
rect 1383 93 1447 157
<< viali >>
rect 1390 100 1440 150
<< locali >>
rect 0 9850 1540 9900
<< locali >>
rect 0 0 1540 50
<< m1 >>
rect 0 50 50 9850
<< m1 >>
rect 1490 50 1540 9850
<< locali >>
rect -7 9843 57 9907
<< m1 >>
rect -7 9843 57 9907
<< viali >>
rect 0 9850 50 9900
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1483 9843 1547 9907
<< m1 >>
rect 1483 9843 1547 9907
<< viali >>
rect 1490 9850 1540 9900
<< locali >>
rect 1483 -7 1547 57
<< m1 >>
rect 1483 -7 1547 57
<< viali >>
rect 1490 0 1540 50
<< locali >>
rect 252 9300 540 9340
<< locali >>
rect 0 9472 1540 9568
<< locali >>
rect -7 9465 57 9575
<< m1 >>
rect -7 9465 57 9575
<< viali >>
rect 0 9472 50 9568
<< locali >>
rect 1483 9465 1547 9575
<< m1 >>
rect 1483 9465 1547 9575
<< viali >>
rect 1490 9472 1540 9568
<< locali >>
rect 0 8832 1540 8928
<< locali >>
rect -7 8825 57 8935
<< m1 >>
rect -7 8825 57 8935
<< viali >>
rect 0 8832 50 8928
<< locali >>
rect 1483 8825 1547 8935
<< m1 >>
rect 1483 8825 1547 8935
<< viali >>
rect 1490 8832 1540 8928
use OTA U2_OTA 
transform 1 0 1590 0 1 0
box 0 0 2886 11510
use temp_affected_current U1_temp_affected_current 
transform 1 0 10316 0 1 0
box 0 0 8726 9970
<< labels >>
flabel locali s 100 9750 1440 9800 0 FreeSans 400 0 0 0 VDD
port 7 nsew signal bidirectional
flabel locali s 0 9850 1540 9900 0 FreeSans 400 0 0 0 VSS
port 8 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1743170539
<< checkpaint >>
rect 0 0 0 0
<< labels >>
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1747235371
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0  diff1_MP3<3> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<2> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 2004
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<1> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 1604
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  diff1_MP3<1>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 1364
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP3<0> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 1604
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  diff1_MP3<0>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 1364
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP4<3> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 2804
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<2> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 2804
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<1> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<0> ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror1_MP2 ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mirror1_MP2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 3604
box 0 0 576 240
use JNWATR_PCH_4C5F0  mirror1_MP1 ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mirror1_MP1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 3604
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN1 ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 292 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN2 ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 904
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1747235371
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWTR_RPPO16  bias1_RH1 ../JNW_TR_SKY130A
timestamp 1747235371
transform 1 0 1644 0 1 200
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH2 ../JNW_TR_SKY130A
timestamp 1747235371
transform 1 0 1644 0 1 3740
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH3 ../JNW_TR_SKY130A
timestamp 1747235371
transform 1 0 1644 0 1 1970
box 0 0 2236 1720
<< m2 >>
rect 820 2187 963 2217
<< m3 >>
rect 820 1787 850 2217
<< m2 >>
rect 820 1787 978 1817
<< m2 >>
rect 372 1787 978 1817
<< m2 >>
rect 244 1787 402 1817
<< m3 >>
rect 244 1787 274 2217
<< m2 >>
rect 244 2187 387 2217
<< m2 >>
rect 813 2180 857 2224
<< m3 >>
rect 813 2180 857 2224
<< via2 >>
rect 820 2187 850 2217
<< m2 >>
rect 813 1780 857 1824
<< m3 >>
rect 813 1780 857 1824
<< via2 >>
rect 820 1787 850 1817
<< m2 >>
rect 237 1780 281 1824
<< m3 >>
rect 237 1780 281 1824
<< via2 >>
rect 244 1787 274 1817
<< m2 >>
rect 237 2180 281 2224
<< m3 >>
rect 237 2180 281 2224
<< via2 >>
rect 244 2187 274 2217
<< m2 >>
rect 820 2987 963 3017
<< m3 >>
rect 820 2587 850 3017
<< m2 >>
rect 820 2587 978 2617
<< m2 >>
rect 372 2587 978 2617
<< m2 >>
rect 244 2587 402 2617
<< m3 >>
rect 244 2587 274 3017
<< m2 >>
rect 244 2987 387 3017
<< m2 >>
rect 813 2980 857 3024
<< m3 >>
rect 813 2980 857 3024
<< via2 >>
rect 820 2987 850 3017
<< m2 >>
rect 813 2580 857 2624
<< m3 >>
rect 813 2580 857 2624
<< via2 >>
rect 820 2587 850 2617
<< m2 >>
rect 237 2580 281 2624
<< m3 >>
rect 237 2580 281 2624
<< via2 >>
rect 244 2587 274 2617
<< m2 >>
rect 237 2980 281 3024
<< m3 >>
rect 237 2980 281 3024
<< via2 >>
rect 244 2987 274 3017
<< m2 >>
rect 1251 523 1410 553
<< m3 >>
rect 1380 523 1410 2457
<< m2 >>
rect 1236 2427 1410 2457
<< m3 >>
rect 1236 2427 1266 2857
<< m2 >>
rect 660 2827 1266 2857
<< m3 >>
rect 660 2442 690 2857
<< m2 >>
rect 1373 516 1417 560
<< m3 >>
rect 1373 516 1417 560
<< via2 >>
rect 1380 523 1410 553
<< m2 >>
rect 1373 2420 1417 2464
<< m3 >>
rect 1373 2420 1417 2464
<< via2 >>
rect 1380 2427 1410 2457
<< m2 >>
rect 1229 2420 1273 2464
<< m3 >>
rect 1229 2420 1273 2464
<< via2 >>
rect 1236 2427 1266 2457
<< m2 >>
rect 1229 2820 1273 2864
<< m3 >>
rect 1229 2820 1273 2864
<< via2 >>
rect 1236 2827 1266 2857
<< m2 >>
rect 653 2820 697 2864
<< m3 >>
rect 653 2820 697 2864
<< via2 >>
rect 660 2827 690 2857
<< m2 >>
rect 387 684 978 714
<< m2 >>
rect 948 684 1266 714
<< m3 >>
rect 1236 684 1266 1658
<< m3 >>
rect 1236 1628 1266 2058
<< m2 >>
rect 660 2028 1266 2058
<< m3 >>
rect 660 1643 690 2058
<< m2 >>
rect 1229 677 1273 721
<< m3 >>
rect 1229 677 1273 721
<< via2 >>
rect 1236 684 1266 714
<< m2 >>
rect 1229 2021 1273 2065
<< m3 >>
rect 1229 2021 1273 2065
<< via2 >>
rect 1236 2028 1266 2058
<< m2 >>
rect 653 2021 697 2065
<< m3 >>
rect 653 2021 697 2065
<< via2 >>
rect 660 2028 690 2058
<< m2 >>
rect 1252 3221 1411 3251
<< m3 >>
rect 1381 2709 1411 3251
<< m2 >>
rect 1045 2709 1411 2739
<< m2 >>
rect 1045 2709 1411 2739
<< m3 >>
rect 1381 2709 1411 3139
<< m2 >>
rect 1045 3109 1411 3139
<< m2 >>
rect 469 3109 1075 3139
<< m2 >>
rect 149 3109 499 3139
<< m3 >>
rect 149 2709 179 3139
<< m2 >>
rect 149 2709 499 2739
<< m2 >>
rect 149 2709 499 2739
<< m3 >>
rect 149 2309 179 2739
<< m2 >>
rect 149 2309 499 2339
<< m2 >>
rect 149 2309 499 2339
<< m3 >>
rect 149 1909 179 2339
<< m2 >>
rect 149 1909 499 1939
<< m2 >>
rect 469 1909 1075 1939
<< m2 >>
rect 1045 1909 1507 1939
<< m3 >>
rect 1477 1909 1507 2339
<< m2 >>
rect 1060 2309 1507 2339
<< m2 >>
rect 1374 3214 1418 3258
<< m3 >>
rect 1374 3214 1418 3258
<< via2 >>
rect 1381 3221 1411 3251
<< m2 >>
rect 1374 2702 1418 2746
<< m3 >>
rect 1374 2702 1418 2746
<< via2 >>
rect 1381 2709 1411 2739
<< m2 >>
rect 1374 2702 1418 2746
<< m3 >>
rect 1374 2702 1418 2746
<< via2 >>
rect 1381 2709 1411 2739
<< m2 >>
rect 1374 3102 1418 3146
<< m3 >>
rect 1374 3102 1418 3146
<< via2 >>
rect 1381 3109 1411 3139
<< m2 >>
rect 142 3102 186 3146
<< m3 >>
rect 142 3102 186 3146
<< via2 >>
rect 149 3109 179 3139
<< m2 >>
rect 142 2702 186 2746
<< m3 >>
rect 142 2702 186 2746
<< via2 >>
rect 149 2709 179 2739
<< m2 >>
rect 142 2702 186 2746
<< m3 >>
rect 142 2702 186 2746
<< via2 >>
rect 149 2709 179 2739
<< m2 >>
rect 142 2302 186 2346
<< m3 >>
rect 142 2302 186 2346
<< via2 >>
rect 149 2309 179 2339
<< m2 >>
rect 142 2302 186 2346
<< m3 >>
rect 142 2302 186 2346
<< via2 >>
rect 149 2309 179 2339
<< m2 >>
rect 142 1902 186 1946
<< m3 >>
rect 142 1902 186 1946
<< via2 >>
rect 149 1909 179 1939
<< m2 >>
rect 1470 1902 1514 1946
<< m3 >>
rect 1470 1902 1514 1946
<< via2 >>
rect 1477 1909 1507 1939
<< m2 >>
rect 1470 2302 1514 2346
<< m3 >>
rect 1470 2302 1514 2346
<< via2 >>
rect 1477 2309 1507 2339
<< m3 >>
rect 3604 1721 3634 3032
<< m2 >>
rect 1620 3002 3634 3032
<< m3 >>
rect 1620 3002 1650 3416
<< m2 >>
rect 948 3386 1650 3416
<< m2 >>
rect 387 3386 978 3416
<< m2 >>
rect 3597 2995 3641 3039
<< m3 >>
rect 3597 2995 3641 3039
<< via2 >>
rect 3604 3002 3634 3032
<< m2 >>
rect 1613 2995 1657 3039
<< m3 >>
rect 1613 2995 1657 3039
<< via2 >>
rect 1620 3002 1650 3032
<< m2 >>
rect 1613 3379 1657 3423
<< m3 >>
rect 1613 3379 1657 3423
<< via2 >>
rect 1620 3386 1650 3416
<< m2 >>
rect 1893 1703 3460 1733
<< m3 >>
rect 3430 1703 3460 5269
<< m2 >>
rect 3430 5239 3621 5269
<< m2 >>
rect 3423 1696 3467 1740
<< m3 >>
rect 3423 1696 3467 1740
<< via2 >>
rect 3430 1703 3460 1733
<< m2 >>
rect 3423 5232 3467 5276
<< m3 >>
rect 3423 5232 3467 5276
<< via2 >>
rect 3430 5239 3460 5269
<< m3 >>
rect 1878 3689 1908 5256
<< m2 >>
rect 1878 3689 3636 3719
<< m3 >>
rect 3606 3480 3636 3719
<< m2 >>
rect 1871 3682 1915 3726
<< m3 >>
rect 1871 3682 1915 3726
<< via2 >>
rect 1878 3689 1908 3719
<< m2 >>
rect 3599 3682 3643 3726
<< m3 >>
rect 3599 3682 3643 3726
<< via2 >>
rect 3606 3689 3636 3719
<< locali >>
rect 100 5510 3980 5560
<< locali >>
rect 100 100 3980 150
<< m1 >>
rect 100 150 150 5510
<< m1 >>
rect 3930 150 3980 5510
<< locali >>
rect 93 5503 157 5567
<< m1 >>
rect 93 5503 157 5567
<< viali >>
rect 100 5510 150 5560
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 3923 5503 3987 5567
<< m1 >>
rect 3923 5503 3987 5567
<< viali >>
rect 3930 5510 3980 5560
<< locali >>
rect 3923 93 3987 157
<< m1 >>
rect 3923 93 3987 157
<< viali >>
rect 3930 100 3980 150
<< locali >>
rect 0 5610 4080 5660
<< locali >>
rect 0 0 4080 50
<< m1 >>
rect 0 50 50 5610
<< m1 >>
rect 4030 50 4080 5610
<< locali >>
rect -7 5603 57 5667
<< m1 >>
rect -7 5603 57 5667
<< viali >>
rect 0 5610 50 5660
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 4023 5603 4087 5667
<< m1 >>
rect 4023 5603 4087 5667
<< viali >>
rect 4030 5610 4080 5660
<< locali >>
rect 4023 -7 4087 57
<< m1 >>
rect 4023 -7 4087 57
<< viali >>
rect 4030 0 4080 50
<< locali >>
rect 1652 3430 1970 3550
<< locali >>
rect 1644 1864 3980 1920
<< locali >>
rect 3923 1857 3987 1927
<< m1 >>
rect 3923 1857 3987 1927
<< viali >>
rect 3930 1864 3980 1920
<< locali >>
rect 1644 200 3980 256
<< locali >>
rect 3923 193 3987 263
<< m1 >>
rect 3923 193 3987 263
<< viali >>
rect 3930 200 3980 256
<< locali >>
rect 1644 5404 3980 5460
<< locali >>
rect 3923 5397 3987 5467
<< m1 >>
rect 3923 5397 3987 5467
<< viali >>
rect 3930 5404 3980 5460
<< locali >>
rect 1644 3740 3980 3796
<< locali >>
rect 3923 3733 3987 3803
<< m1 >>
rect 3923 3733 3987 3803
<< viali >>
rect 3930 3740 3980 3796
<< locali >>
rect 1644 3634 3980 3690
<< locali >>
rect 3923 3627 3987 3697
<< m1 >>
rect 3923 3627 3987 3697
<< viali >>
rect 3930 3634 3980 3690
<< locali >>
rect 1644 1970 3980 2026
<< locali >>
rect 3923 1963 3987 2033
<< m1 >>
rect 3923 1963 3987 2033
<< viali >>
rect 3930 1970 3980 2026
<< locali >>
rect 820 3504 1108 3544
<< locali >>
rect 244 3504 532 3544
<< locali >>
rect 628 3384 788 3424
<< locali >>
rect 244 804 532 844
<< locali >>
rect 628 684 788 724
<< locali >>
rect 820 804 1108 844
<< locali >>
rect 0 1436 1352 1532
<< locali >>
rect -7 1429 57 1539
<< m1 >>
rect -7 1429 57 1539
<< viali >>
rect 0 1436 50 1532
<< locali >>
rect 0 3676 1352 3772
<< locali >>
rect -7 3669 57 3779
<< m1 >>
rect -7 3669 57 3779
<< viali >>
rect 0 3676 50 3772
<< locali >>
rect 100 976 1352 1072
<< locali >>
rect 93 969 157 1079
<< m1 >>
rect 93 969 157 1079
<< viali >>
rect 100 976 150 1072
<< locali >>
rect 100 336 1352 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< m1 >>
rect 365 2177 411 2231
<< m2 >>
rect 365 2177 411 2231
<< via1 >>
rect 372 2184 404 2224
<< m1 >>
rect 941 2177 987 2231
<< m2 >>
rect 941 2177 987 2231
<< via1 >>
rect 948 2184 980 2224
<< m1 >>
rect 365 1777 411 1831
<< m2 >>
rect 365 1777 411 1831
<< via1 >>
rect 372 1784 404 1824
<< m1 >>
rect 365 1777 411 1831
<< m2 >>
rect 365 1777 411 1831
<< via1 >>
rect 372 1784 404 1824
<< m1 >>
rect 941 1777 987 1831
<< m2 >>
rect 941 1777 987 1831
<< via1 >>
rect 948 1784 980 1824
<< m1 >>
rect 941 1777 987 1831
<< m2 >>
rect 941 1777 987 1831
<< via1 >>
rect 948 1784 980 1824
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 941 2977 987 3031
<< m2 >>
rect 941 2977 987 3031
<< via1 >>
rect 948 2984 980 3024
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< m3 >>
rect 621 2817 731 2871
<< via2 >>
rect 628 2824 724 2864
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< m3 >>
rect 1197 2817 1307 2871
<< via2 >>
rect 1204 2824 1300 2864
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 1197 2417 1307 2471
<< m2 >>
rect 1197 2417 1307 2471
<< m3 >>
rect 1197 2417 1307 2471
<< via2 >>
rect 1204 2424 1300 2464
<< via1 >>
rect 1204 2424 1300 2464
<< m1 >>
rect 621 2417 731 2471
<< m2 >>
rect 621 2417 731 2471
<< m3 >>
rect 621 2417 731 2471
<< via2 >>
rect 628 2424 724 2464
<< via1 >>
rect 628 2424 724 2464
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 621 2017 731 2071
<< m2 >>
rect 621 2017 731 2071
<< m3 >>
rect 621 2017 731 2071
<< via2 >>
rect 628 2024 724 2064
<< via1 >>
rect 628 2024 724 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< m3 >>
rect 1197 2017 1307 2071
<< via2 >>
rect 1204 2024 1300 2064
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 1197 2017 1307 2071
<< m2 >>
rect 1197 2017 1307 2071
<< via1 >>
rect 1204 2024 1300 2064
<< m1 >>
rect 621 1617 731 1671
<< m2 >>
rect 621 1617 731 1671
<< m3 >>
rect 621 1617 731 1671
<< via2 >>
rect 628 1624 724 1664
<< via1 >>
rect 628 1624 724 1664
<< m1 >>
rect 1197 1617 1307 1671
<< m2 >>
rect 1197 1617 1307 1671
<< m3 >>
rect 1197 1617 1307 1671
<< via2 >>
rect 1204 1624 1300 1664
<< via1 >>
rect 1204 1624 1300 1664
<< m1 >>
rect 1197 1617 1307 1671
<< m2 >>
rect 1197 1617 1307 1671
<< m3 >>
rect 1197 1617 1307 1671
<< via2 >>
rect 1204 1624 1300 1664
<< via1 >>
rect 1204 1624 1300 1664
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 429 2297 539 2351
<< m2 >>
rect 429 2297 539 2351
<< via1 >>
rect 436 2304 532 2344
<< m1 >>
rect 1005 2297 1115 2351
<< m2 >>
rect 1005 2297 1115 2351
<< via1 >>
rect 1012 2304 1108 2344
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 429 1897 539 1951
<< m2 >>
rect 429 1897 539 1951
<< via1 >>
rect 436 1904 532 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 1005 1897 1115 1951
<< m2 >>
rect 1005 1897 1115 1951
<< via1 >>
rect 1012 1904 1108 1944
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 429 3097 539 3151
<< m2 >>
rect 429 3097 539 3151
<< via1 >>
rect 436 3104 532 3144
<< m1 >>
rect 1005 3097 1115 3151
<< m2 >>
rect 1005 3097 1115 3151
<< via1 >>
rect 1012 3104 1108 3144
<< m1 >>
rect 1005 3097 1115 3151
<< m2 >>
rect 1005 3097 1115 3151
<< via1 >>
rect 1012 3104 1108 3144
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 1005 2697 1115 2751
<< m2 >>
rect 1005 2697 1115 2751
<< via1 >>
rect 1012 2704 1108 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 429 2697 539 2751
<< m2 >>
rect 429 2697 539 2751
<< via1 >>
rect 436 2704 532 2744
<< m1 >>
rect 1197 3217 1307 3271
<< m2 >>
rect 1197 3217 1307 3271
<< via1 >>
rect 1204 3224 1300 3264
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 365 3377 411 3431
<< m2 >>
rect 365 3377 411 3431
<< via1 >>
rect 372 3384 404 3424
<< locali >>
rect 3547 1653 3705 1787
<< m1 >>
rect 3547 1653 3705 1787
<< m2 >>
rect 3547 1653 3705 1787
<< m3 >>
rect 3547 1653 3705 1787
<< via2 >>
rect 3554 1660 3698 1780
<< via1 >>
rect 3554 1660 3698 1780
<< viali >>
rect 3554 1660 3698 1780
<< locali >>
rect 1819 1653 1977 1787
<< m1 >>
rect 1819 1653 1977 1787
<< m2 >>
rect 1819 1653 1977 1787
<< via1 >>
rect 1826 1660 1970 1780
<< viali >>
rect 1826 1660 1970 1780
<< locali >>
rect 3547 5193 3705 5327
<< m1 >>
rect 3547 5193 3705 5327
<< m2 >>
rect 3547 5193 3705 5327
<< via1 >>
rect 3554 5200 3698 5320
<< viali >>
rect 3554 5200 3698 5320
<< locali >>
rect 1819 5193 1977 5327
<< m1 >>
rect 1819 5193 1977 5327
<< m2 >>
rect 1819 5193 1977 5327
<< m3 >>
rect 1819 5193 1977 5327
<< via2 >>
rect 1826 5200 1970 5320
<< via1 >>
rect 1826 5200 1970 5320
<< viali >>
rect 1826 5200 1970 5320
<< locali >>
rect 3547 3423 3705 3557
<< m1 >>
rect 3547 3423 3705 3557
<< m2 >>
rect 3547 3423 3705 3557
<< m3 >>
rect 3547 3423 3705 3557
<< via2 >>
rect 3554 3430 3698 3550
<< via1 >>
rect 3554 3430 3698 3550
<< viali >>
rect 3554 3430 3698 3550
<< labels >>
flabel m2 s 820 2187 963 2217 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 820 2987 963 3017 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 0 5610 4080 5660 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 100 5510 3980 5560 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m2 s 1251 523 1410 553 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1729505989
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 x1 ../JNW_ATR_SKY130A
transform 0 -1 400 1 0 9856
box 0 0 832 400
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform -1 0 512 0 -1 9024
box 0 0 512 400
use JNWTR_CAPX1 x4 ../JNW_TR_SKY130A
transform -1 0 2332 0 -1 8048
box 0 0 540 540
use JNWTR_RES2 x3 ../JNW_TR_SKY130A
transform 0 -1 3112 1 0 8624
box 0 0 324 1320
use JNWATR_NCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 0 -1 992 1 0 10000
box 0 0 576 400
use JNWATR_NCH_4C5F0 x3 ../JNW_ATR_SKY130A
transform 0 -1 912 1 0 9240
box 0 0 576 400
use JNWATR_PCH_4C5F0 x7 ../JNW_ATR_SKY130A
transform -1 0 2064 0 -1 9024
box 0 0 576 400
use JNWATR_PCH_4C5F0 x9 ../JNW_ATR_SKY130A
transform -1 0 1488 0 -1 9024
box 0 0 576 400
use JNWATR_PCH_4C5F0 x8 ../JNW_ATR_SKY130A
transform -1 0 2064 0 -1 9424
box 0 0 576 400
use JNWATR_PCH_4C5F0 x5 ../JNW_ATR_SKY130A
transform 0 1 1792 -1 0 10000
box 0 0 576 400
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform 0 1 688 -1 0 8624
box 0 0 576 400
use JNWATR_NCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 512 0 1 512
box 0 0 576 400
use JNWATR_NCH_4C5F0 x10 ../JNW_ATR_SKY130A
transform 0 -1 1488 1 0 8624
box 0 0 576 400
use JNWATR_NCH_4C5F0 x11 ../JNW_ATR_SKY130A
transform 0 1 1088 -1 0 8624
box 0 0 576 400
use JNWATR_PCH_4C5F0 x12 ../JNW_ATR_SKY130A
transform 0 1 1392 -1 0 10000
box 0 0 576 400
use JNWATR_PCH_4C5F0 x13 ../JNW_ATR_SKY130A
transform -1 0 1488 0 -1 9424
box 0 0 576 400
<< labels >>
<< properties >>
<< end >>
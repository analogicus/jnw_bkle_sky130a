magic
tech sky130A
magscale 1 1
timestamp 1737716231
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 MN7 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN8 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP5 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 900
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP6 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 900
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 100
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP2 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 100
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN10 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN9 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN11 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 2100
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN12 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 2100
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP3 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 500
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP4 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 500
box 0 0 576 400
<< m1 >>
rect 1637 1793 1747 1847
<< m2 >>
rect 1637 1793 1747 1847
<< m3 >>
rect 1637 1793 1747 1847
<< via2 >>
rect 1644 1800 1740 1840
<< via1 >>
rect 1644 1800 1740 1840
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< m3 >>
rect 1061 1793 1171 1847
<< via2 >>
rect 1068 1800 1164 1840
<< via1 >>
rect 1068 1800 1164 1840
<< locali >>
rect 869 1673 979 1727
<< m1 >>
rect 869 1673 979 1727
<< m2 >>
rect 869 1673 979 1727
<< via1 >>
rect 876 1680 972 1720
<< viali >>
rect 876 1680 972 1720
<< m1 >>
rect 997 1073 1043 1127
<< m2 >>
rect 997 1073 1043 1127
<< via1 >>
rect 1004 1080 1036 1120
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< m3 >>
rect 1253 913 1363 967
<< via2 >>
rect 1260 920 1356 960
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< locali >>
rect 869 1073 979 1127
<< m1 >>
rect 869 1073 979 1127
<< m2 >>
rect 869 1073 979 1127
<< via1 >>
rect 876 1080 972 1120
<< viali >>
rect 876 1080 972 1120
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< m3 >>
rect 1637 393 1747 447
<< via2 >>
rect 1644 400 1740 440
<< via1 >>
rect 1644 400 1740 440
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 997 273 1043 327
<< m2 >>
rect 997 273 1043 327
<< via1 >>
rect 1004 280 1036 320
<< m1 >>
rect 1253 113 1363 167
<< m2 >>
rect 1253 113 1363 167
<< m3 >>
rect 1253 113 1363 167
<< via2 >>
rect 1260 120 1356 160
<< via1 >>
rect 1260 120 1356 160
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< m3 >>
rect 1061 393 1171 447
<< via2 >>
rect 1068 400 1164 440
<< via1 >>
rect 1068 400 1164 440
<< locali >>
rect 869 273 979 327
<< m1 >>
rect 869 273 979 327
<< m2 >>
rect 869 273 979 327
<< via1 >>
rect 876 280 972 320
<< viali >>
rect 876 280 972 320
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< m3 >>
rect 1061 2793 1171 2847
<< via2 >>
rect 1068 2800 1164 2840
<< via1 >>
rect 1068 2800 1164 2840
<< locali >>
rect 869 2673 979 2727
<< m1 >>
rect 869 2673 979 2727
<< m2 >>
rect 869 2673 979 2727
<< via1 >>
rect 876 2680 972 2720
<< viali >>
rect 876 2680 972 2720
<< m1 >>
rect 1573 2673 1619 2727
<< m2 >>
rect 1573 2673 1619 2727
<< via1 >>
rect 1580 2680 1612 2720
<< m1 >>
rect 1829 2513 1939 2567
<< m2 >>
rect 1829 2513 1939 2567
<< m3 >>
rect 1829 2513 1939 2567
<< via2 >>
rect 1836 2520 1932 2560
<< via1 >>
rect 1836 2520 1932 2560
<< m1 >>
rect 1637 2793 1747 2847
<< m2 >>
rect 1637 2793 1747 2847
<< m3 >>
rect 1637 2793 1747 2847
<< via2 >>
rect 1644 2800 1740 2840
<< via1 >>
rect 1644 2800 1740 2840
<< locali >>
rect 1445 2673 1555 2727
<< m1 >>
rect 1445 2673 1555 2727
<< m2 >>
rect 1445 2673 1555 2727
<< via1 >>
rect 1452 2680 1548 2720
<< viali >>
rect 1452 2680 1548 2720
<< m1 >>
rect 997 2273 1043 2327
<< m2 >>
rect 997 2273 1043 2327
<< via1 >>
rect 1004 2280 1036 2320
<< m1 >>
rect 1253 2113 1363 2167
<< m2 >>
rect 1253 2113 1363 2167
<< m3 >>
rect 1253 2113 1363 2167
<< via2 >>
rect 1260 2120 1356 2160
<< via1 >>
rect 1260 2120 1356 2160
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< locali >>
rect 869 2273 979 2327
<< m1 >>
rect 869 2273 979 2327
<< m2 >>
rect 869 2273 979 2327
<< via1 >>
rect 876 2280 972 2320
<< viali >>
rect 876 2280 972 2320
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< m3 >>
rect 1637 2393 1747 2447
<< via2 >>
rect 1644 2400 1740 2440
<< via1 >>
rect 1644 2400 1740 2440
<< locali >>
rect 1445 2273 1555 2327
<< m1 >>
rect 1445 2273 1555 2327
<< m2 >>
rect 1445 2273 1555 2327
<< via1 >>
rect 1452 2280 1548 2320
<< viali >>
rect 1452 2280 1548 2320
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< locali >>
rect 869 673 979 727
<< m1 >>
rect 869 673 979 727
<< m2 >>
rect 869 673 979 727
<< via1 >>
rect 876 680 972 720
<< viali >>
rect 876 680 972 720
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< m3 >>
rect 1445 1673 1555 1727
<< via2 >>
rect 1452 1680 1548 1720
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1637 1793 1747 1847
<< m2 >>
rect 1637 1793 1747 1847
<< via1 >>
rect 1644 1800 1740 1840
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< m3 >>
rect 1445 1673 1555 1727
<< via2 >>
rect 1452 1680 1548 1720
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1253 113 1363 167
<< m2 >>
rect 1253 113 1363 167
<< via1 >>
rect 1260 120 1356 160
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< m3 >>
rect 1253 513 1363 567
<< via2 >>
rect 1260 520 1356 560
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< m3 >>
rect 1445 1673 1555 1727
<< via2 >>
rect 1452 1680 1548 1720
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1637 1793 1747 1847
<< m2 >>
rect 1637 1793 1747 1847
<< via1 >>
rect 1644 1800 1740 1840
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< m3 >>
rect 1445 1673 1555 1727
<< via2 >>
rect 1452 1680 1548 1720
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< m3 >>
rect 1445 1673 1555 1727
<< via2 >>
rect 1452 1680 1548 1720
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< m3 >>
rect 1061 1793 1171 1847
<< via2 >>
rect 1068 1800 1164 1840
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< m3 >>
rect 1253 913 1363 967
<< via2 >>
rect 1260 920 1356 960
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< m3 >>
rect 1061 1793 1171 1847
<< via2 >>
rect 1068 1800 1164 1840
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< via1 >>
rect 1068 1800 1164 1840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< m3 >>
rect 1637 393 1747 447
<< via2 >>
rect 1644 400 1740 440
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< m3 >>
rect 1061 393 1171 447
<< via2 >>
rect 1068 400 1164 440
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< m3 >>
rect 1253 913 1363 967
<< via2 >>
rect 1260 920 1356 960
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< m3 >>
rect 1445 1073 1555 1127
<< via2 >>
rect 1452 1080 1548 1120
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< m3 >>
rect 1445 1073 1555 1127
<< via2 >>
rect 1452 1080 1548 1120
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< m3 >>
rect 1445 273 1555 327
<< via2 >>
rect 1452 280 1548 320
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 1253 113 1363 167
<< m2 >>
rect 1253 113 1363 167
<< via1 >>
rect 1260 120 1356 160
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< m3 >>
rect 1445 273 1555 327
<< via2 >>
rect 1452 280 1548 320
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< m3 >>
rect 1253 1513 1363 1567
<< via2 >>
rect 1260 1520 1356 1560
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< via1 >>
rect 1260 920 1356 960
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< m3 >>
rect 1445 273 1555 327
<< via2 >>
rect 1452 280 1548 320
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 1253 2113 1363 2167
<< m2 >>
rect 1253 2113 1363 2167
<< via1 >>
rect 1260 2120 1356 2160
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 2273 1555 2327
<< m1 >>
rect 1445 2273 1555 2327
<< m2 >>
rect 1445 2273 1555 2327
<< via1 >>
rect 1452 2280 1548 2320
<< viali >>
rect 1452 2280 1548 2320
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< m3 >>
rect 1445 273 1555 327
<< via2 >>
rect 1452 280 1548 320
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1253 113 1363 167
<< m2 >>
rect 1253 113 1363 167
<< via1 >>
rect 1260 120 1356 160
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< m3 >>
rect 1253 513 1363 567
<< via2 >>
rect 1260 520 1356 560
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< via1 >>
rect 1068 400 1164 440
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 997 273 1043 327
<< m2 >>
rect 997 273 1043 327
<< via1 >>
rect 1004 280 1036 320
<< m1 >>
rect 997 673 1043 727
<< m2 >>
rect 997 673 1043 727
<< via1 >>
rect 1004 680 1036 720
<< m1 >>
rect 997 673 1043 727
<< m2 >>
rect 997 673 1043 727
<< m3 >>
rect 997 673 1043 727
<< via2 >>
rect 1004 680 1036 720
<< via1 >>
rect 1004 680 1036 720
<< m1 >>
rect 997 673 1043 727
<< m2 >>
rect 997 673 1043 727
<< via1 >>
rect 1004 680 1036 720
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1253 2513 1363 2567
<< m2 >>
rect 1253 2513 1363 2567
<< m3 >>
rect 1253 2513 1363 2567
<< via2 >>
rect 1260 2520 1356 2560
<< via1 >>
rect 1260 2520 1356 2560
<< m1 >>
rect 1829 2513 1939 2567
<< m2 >>
rect 1829 2513 1939 2567
<< m3 >>
rect 1829 2513 1939 2567
<< via2 >>
rect 1836 2520 1932 2560
<< via1 >>
rect 1836 2520 1932 2560
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< m3 >>
rect 1061 2793 1171 2847
<< via2 >>
rect 1068 2800 1164 2840
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1637 2793 1747 2847
<< m2 >>
rect 1637 2793 1747 2847
<< m3 >>
rect 1637 2793 1747 2847
<< via2 >>
rect 1644 2800 1740 2840
<< via1 >>
rect 1644 2800 1740 2840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< m3 >>
rect 1061 2793 1171 2847
<< via2 >>
rect 1068 2800 1164 2840
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2793 1171 2847
<< m2 >>
rect 1061 2793 1171 2847
<< via1 >>
rect 1068 2800 1164 2840
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< m3 >>
rect 1637 2393 1747 2447
<< via2 >>
rect 1644 2400 1740 2440
<< via1 >>
rect 1644 2400 1740 2440
<< locali >>
rect 1445 2673 1555 2727
<< m1 >>
rect 1445 2673 1555 2727
<< m2 >>
rect 1445 2673 1555 2727
<< m3 >>
rect 1445 2673 1555 2727
<< via2 >>
rect 1452 2680 1548 2720
<< via1 >>
rect 1452 2680 1548 2720
<< viali >>
rect 1452 2680 1548 2720
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1637 2793 1747 2847
<< m2 >>
rect 1637 2793 1747 2847
<< via1 >>
rect 1644 2800 1740 2840
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< via1 >>
rect 1644 2400 1740 2440
<< m1 >>
rect 1253 2113 1363 2167
<< m2 >>
rect 1253 2113 1363 2167
<< via1 >>
rect 1260 2120 1356 2160
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< m3 >>
rect 1637 2393 1747 2447
<< via2 >>
rect 1644 2400 1740 2440
<< via1 >>
rect 1644 2400 1740 2440
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< via1 >>
rect 1644 2400 1740 2440
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< m3 >>
rect 1637 2393 1747 2447
<< via2 >>
rect 1644 2400 1740 2440
<< via1 >>
rect 1644 2400 1740 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1061 2393 1171 2447
<< m2 >>
rect 1061 2393 1171 2447
<< m3 >>
rect 1061 2393 1171 2447
<< via2 >>
rect 1068 2400 1164 2440
<< via1 >>
rect 1068 2400 1164 2440
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< m3 >>
rect 1637 2393 1747 2447
<< via2 >>
rect 1644 2400 1740 2440
<< via1 >>
rect 1644 2400 1740 2440
<< m1 >>
rect 1637 2393 1747 2447
<< m2 >>
rect 1637 2393 1747 2447
<< via1 >>
rect 1644 2400 1740 2440
<< m3 >>
rect 1485 1805 1692 1835
<< m2 >>
rect 1485 1700 1515 1835
<< m2 >>
rect 1478 1798 1522 1842
<< m3 >>
rect 1478 1798 1522 1842
<< via2 >>
rect 1485 1805 1515 1835
<< m3 >>
rect 909 1805 1116 1835
<< m2 >>
rect 909 1700 939 1835
<< m2 >>
rect 902 1798 946 1842
<< m3 >>
rect 902 1798 946 1842
<< via2 >>
rect 909 1805 939 1835
<< m3 >>
rect 1005 925 1308 955
<< m2 >>
rect 1005 925 1035 1100
<< m2 >>
rect 998 918 1042 962
<< m3 >>
rect 998 918 1042 962
<< via2 >>
rect 1005 925 1035 955
<< m3 >>
rect 909 1205 1116 1235
<< m2 >>
rect 909 1100 939 1235
<< m2 >>
rect 902 1198 946 1242
<< m3 >>
rect 902 1198 946 1242
<< via2 >>
rect 909 1205 939 1235
<< m3 >>
rect 1485 1205 1692 1235
<< m2 >>
rect 1485 1100 1515 1235
<< m2 >>
rect 1478 1198 1522 1242
<< m3 >>
rect 1478 1198 1522 1242
<< via2 >>
rect 1485 1205 1515 1235
<< m3 >>
rect 1485 405 1692 435
<< m2 >>
rect 1485 300 1515 435
<< m2 >>
rect 1478 398 1522 442
<< m3 >>
rect 1478 398 1522 442
<< via2 >>
rect 1485 405 1515 435
<< m3 >>
rect 1005 125 1308 155
<< m2 >>
rect 1005 125 1035 300
<< m2 >>
rect 998 118 1042 162
<< m3 >>
rect 998 118 1042 162
<< via2 >>
rect 1005 125 1035 155
<< m3 >>
rect 909 405 1116 435
<< m2 >>
rect 909 300 939 435
<< m2 >>
rect 902 398 946 442
<< m3 >>
rect 902 398 946 442
<< via2 >>
rect 909 405 939 435
<< m3 >>
rect 909 2805 1116 2835
<< m2 >>
rect 909 2700 939 2835
<< m2 >>
rect 902 2798 946 2842
<< m3 >>
rect 902 2798 946 2842
<< via2 >>
rect 909 2805 939 2835
<< m3 >>
rect 1581 2525 1884 2555
<< m2 >>
rect 1581 2525 1611 2700
<< m2 >>
rect 1574 2518 1618 2562
<< m3 >>
rect 1574 2518 1618 2562
<< via2 >>
rect 1581 2525 1611 2555
<< m3 >>
rect 1485 2805 1692 2835
<< m2 >>
rect 1485 2700 1515 2835
<< m2 >>
rect 1478 2798 1522 2842
<< m3 >>
rect 1478 2798 1522 2842
<< via2 >>
rect 1485 2805 1515 2835
<< m3 >>
rect 1005 2125 1308 2155
<< m2 >>
rect 1005 2125 1035 2300
<< m2 >>
rect 998 2118 1042 2162
<< m3 >>
rect 998 2118 1042 2162
<< via2 >>
rect 1005 2125 1035 2155
<< m3 >>
rect 909 2405 1116 2435
<< m2 >>
rect 909 2300 939 2435
<< m2 >>
rect 902 2398 946 2442
<< m3 >>
rect 902 2398 946 2442
<< via2 >>
rect 909 2405 939 2435
<< m3 >>
rect 1485 2405 1692 2435
<< m2 >>
rect 1485 2300 1515 2435
<< m2 >>
rect 1478 2398 1522 2442
<< m3 >>
rect 1478 2398 1522 2442
<< via2 >>
rect 1485 2405 1515 2435
<< m3 >>
rect 1485 805 1692 835
<< m2 >>
rect 1485 700 1515 835
<< m2 >>
rect 1478 798 1522 842
<< m3 >>
rect 1478 798 1522 842
<< via2 >>
rect 1485 805 1515 835
<< m3 >>
rect 909 805 1116 835
<< m2 >>
rect 909 700 939 835
<< m2 >>
rect 902 798 946 842
<< m3 >>
rect 902 798 946 842
<< via2 >>
rect 909 805 939 835
<< m3 >>
rect 1101 1685 1500 1715
<< m2 >>
rect 1101 1685 1131 1820
<< m2 >>
rect 1094 1678 1138 1722
<< m3 >>
rect 1094 1678 1138 1722
<< via2 >>
rect 1101 1685 1131 1715
<< m2 >>
rect 1677 1206 1707 1820
<< m2 >>
rect 1677 1206 1707 1236
<< m2 >>
rect 1677 405 1707 1236
<< m2 >>
rect 1677 405 1707 420
<< m2 >>
rect 1485 1684 1515 1700
<< m3 >>
rect 1294 1684 1515 1714
<< m2 >>
rect 1294 524 1324 1714
<< m3 >>
rect 1293 524 1324 554
<< m2 >>
rect 1293 140 1323 554
<< m2 >>
rect 1478 1677 1522 1707
<< m3 >>
rect 1478 1677 1522 1707
<< via2 >>
rect 1485 1684 1515 1700
<< m2 >>
rect 1287 1677 1331 1721
<< m3 >>
rect 1287 1677 1331 1721
<< via2 >>
rect 1294 1684 1324 1714
<< m2 >>
rect 1287 517 1331 561
<< m3 >>
rect 1287 517 1331 561
<< via2 >>
rect 1294 524 1324 554
<< m2 >>
rect 1286 517 1330 561
<< m3 >>
rect 1286 517 1330 561
<< via2 >>
rect 1293 524 1323 554
<< m3 >>
rect 1102 1685 1500 1715
<< m2 >>
rect 1102 1685 1132 2436
<< m3 >>
rect 1101 2406 1132 2436
<< m2 >>
rect 1101 2406 1131 2820
<< m2 >>
rect 1095 1678 1139 1722
<< m3 >>
rect 1095 1678 1139 1722
<< via2 >>
rect 1102 1685 1132 1715
<< m2 >>
rect 1095 2399 1139 2443
<< m3 >>
rect 1095 2399 1139 2443
<< via2 >>
rect 1102 2406 1132 2436
<< m2 >>
rect 1094 2399 1138 2443
<< m3 >>
rect 1094 2399 1138 2443
<< via2 >>
rect 1101 2406 1131 2436
<< m2 >>
rect 1677 1207 1707 1820
<< m2 >>
rect 1677 1207 1707 1237
<< m2 >>
rect 1677 1204 1707 1237
<< m2 >>
rect 1677 1204 1707 1234
<< m2 >>
rect 1677 820 1707 1234
<< m3 >>
rect 1483 1685 1500 1715
<< m2 >>
rect 1483 1684 1513 1715
<< m3 >>
rect 1295 1684 1513 1714
<< m2 >>
rect 1295 1683 1325 1714
<< m3 >>
rect 1102 1683 1325 1713
<< m2 >>
rect 1102 1204 1132 1713
<< m3 >>
rect 1101 1204 1132 1234
<< m2 >>
rect 1101 820 1131 1234
<< m2 >>
rect 1476 1678 1507 1722
<< m3 >>
rect 1476 1678 1507 1722
<< via2 >>
rect 1483 1685 1500 1715
<< m2 >>
rect 1476 1677 1520 1721
<< m3 >>
rect 1476 1677 1520 1721
<< via2 >>
rect 1483 1684 1513 1714
<< m2 >>
rect 1288 1677 1332 1721
<< m3 >>
rect 1288 1677 1332 1721
<< via2 >>
rect 1295 1684 1325 1714
<< m2 >>
rect 1288 1676 1332 1720
<< m3 >>
rect 1288 1676 1332 1720
<< via2 >>
rect 1295 1683 1325 1713
<< m2 >>
rect 1095 1676 1139 1720
<< m3 >>
rect 1095 1676 1139 1720
<< via2 >>
rect 1102 1683 1132 1713
<< m2 >>
rect 1095 1197 1139 1241
<< m3 >>
rect 1095 1197 1139 1241
<< via2 >>
rect 1102 1204 1132 1234
<< m2 >>
rect 1094 1197 1138 1241
<< m3 >>
rect 1094 1197 1138 1241
<< via2 >>
rect 1101 1204 1131 1234
<< m3 >>
rect 1116 1805 1132 1835
<< m2 >>
rect 1102 925 1132 1835
<< m3 >>
rect 1102 925 1308 955
<< m2 >>
rect 1109 1798 1139 1842
<< m3 >>
rect 1109 1798 1139 1842
<< via2 >>
rect 1116 1805 1132 1835
<< m2 >>
rect 1095 918 1139 962
<< m3 >>
rect 1095 918 1139 962
<< via2 >>
rect 1102 925 1132 955
<< m2 >>
rect 1101 1804 1131 1820
<< m3 >>
rect 1101 1804 1131 1834
<< m2 >>
rect 1101 1208 1131 1834
<< m3 >>
rect 1101 1208 1705 1238
<< m2 >>
rect 1675 1205 1705 1238
<< m3 >>
rect 1675 1205 1692 1235
<< m2 >>
rect 1094 1797 1138 1827
<< m3 >>
rect 1094 1797 1138 1827
<< via2 >>
rect 1101 1804 1131 1820
<< m2 >>
rect 1094 1797 1138 1841
<< m3 >>
rect 1094 1797 1138 1841
<< via2 >>
rect 1101 1804 1131 1834
<< m2 >>
rect 1094 1201 1138 1245
<< m3 >>
rect 1094 1201 1138 1245
<< via2 >>
rect 1101 1208 1131 1238
<< m2 >>
rect 1668 1201 1712 1245
<< m3 >>
rect 1668 1201 1712 1245
<< via2 >>
rect 1675 1208 1705 1238
<< m2 >>
rect 1668 1198 1699 1242
<< m3 >>
rect 1668 1198 1699 1242
<< via2 >>
rect 1675 1205 1692 1235
<< m2 >>
rect 1101 1820 1131 2433
<< m2 >>
rect 1101 2403 1131 2433
<< m2 >>
rect 1101 2403 1131 2835
<< m2 >>
rect 1101 2805 1131 2820
<< m2 >>
rect 1101 807 1131 1820
<< m3 >>
rect 1101 807 1705 837
<< m2 >>
rect 1675 805 1705 837
<< m3 >>
rect 1675 805 1707 835
<< m2 >>
rect 1677 820 1707 835
<< m2 >>
rect 1094 800 1138 844
<< m3 >>
rect 1094 800 1138 844
<< via2 >>
rect 1101 807 1131 837
<< m2 >>
rect 1668 800 1712 844
<< m3 >>
rect 1668 800 1712 844
<< via2 >>
rect 1675 807 1705 837
<< m2 >>
rect 1668 798 1712 842
<< m3 >>
rect 1668 798 1712 842
<< via2 >>
rect 1675 805 1705 835
<< m2 >>
rect 1670 813 1714 842
<< m3 >>
rect 1670 813 1714 842
<< via2 >>
rect 1677 820 1707 835
<< m2 >>
rect 1101 807 1131 1820
<< m2 >>
rect 1101 807 1131 837
<< m2 >>
rect 1101 805 1131 837
<< m2 >>
rect 1101 805 1131 820
<< m3 >>
rect 1116 1205 1513 1235
<< m2 >>
rect 1483 1205 1513 1235
<< m3 >>
rect 1483 1205 1515 1235
<< m2 >>
rect 1485 1205 1515 1235
<< m3 >>
rect 1485 1205 1692 1235
<< m2 >>
rect 1476 1198 1520 1242
<< m3 >>
rect 1476 1198 1520 1242
<< via2 >>
rect 1483 1205 1513 1235
<< m2 >>
rect 1476 1198 1520 1242
<< m3 >>
rect 1476 1198 1520 1242
<< via2 >>
rect 1483 1205 1513 1235
<< m2 >>
rect 1478 1198 1522 1242
<< m3 >>
rect 1478 1198 1522 1242
<< via2 >>
rect 1485 1205 1515 1235
<< m2 >>
rect 1478 1198 1522 1242
<< m3 >>
rect 1478 1198 1522 1242
<< via2 >>
rect 1485 1205 1515 1235
<< m3 >>
rect 1116 1205 1132 1235
<< m2 >>
rect 1102 1204 1132 1235
<< m3 >>
rect 1102 1204 1133 1234
<< m2 >>
rect 1103 406 1133 1234
<< m3 >>
rect 1103 406 1707 436
<< m2 >>
rect 1677 420 1707 436
<< m2 >>
rect 1109 1198 1139 1242
<< m3 >>
rect 1109 1198 1139 1242
<< via2 >>
rect 1116 1205 1132 1235
<< m2 >>
rect 1095 1197 1139 1241
<< m3 >>
rect 1095 1197 1139 1241
<< via2 >>
rect 1102 1204 1132 1234
<< m2 >>
rect 1096 1197 1140 1241
<< m3 >>
rect 1096 1197 1140 1241
<< via2 >>
rect 1103 1204 1133 1234
<< m2 >>
rect 1096 399 1140 443
<< m3 >>
rect 1096 399 1140 443
<< via2 >>
rect 1103 406 1133 436
<< m2 >>
rect 1670 413 1714 443
<< m3 >>
rect 1670 413 1714 443
<< via2 >>
rect 1677 420 1707 436
<< m2 >>
rect 1101 1204 1131 1220
<< m2 >>
rect 1101 1204 1131 1234
<< m2 >>
rect 1101 405 1131 1234
<< m2 >>
rect 1101 405 1131 420
<< m2 >>
rect 1293 807 1323 940
<< m3 >>
rect 1293 807 1706 837
<< m2 >>
rect 1676 805 1706 837
<< m3 >>
rect 1676 805 1692 835
<< m2 >>
rect 1286 800 1330 844
<< m3 >>
rect 1286 800 1330 844
<< via2 >>
rect 1293 807 1323 837
<< m2 >>
rect 1669 800 1713 844
<< m3 >>
rect 1669 800 1713 844
<< via2 >>
rect 1676 807 1706 837
<< m2 >>
rect 1669 798 1699 842
<< m3 >>
rect 1669 798 1699 842
<< via2 >>
rect 1676 805 1692 835
<< m3 >>
rect 1116 1205 1134 1235
<< m2 >>
rect 1104 1204 1134 1235
<< m3 >>
rect 1104 1204 1135 1234
<< m2 >>
rect 1105 807 1135 1234
<< m3 >>
rect 1105 807 1516 837
<< m2 >>
rect 1486 805 1516 837
<< m3 >>
rect 1486 805 1692 835
<< m2 >>
rect 1109 1198 1141 1242
<< m3 >>
rect 1109 1198 1141 1242
<< via2 >>
rect 1116 1205 1134 1235
<< m2 >>
rect 1097 1197 1141 1241
<< m3 >>
rect 1097 1197 1141 1241
<< via2 >>
rect 1104 1204 1134 1234
<< m2 >>
rect 1098 1197 1142 1241
<< m3 >>
rect 1098 1197 1142 1241
<< via2 >>
rect 1105 1204 1135 1234
<< m2 >>
rect 1098 800 1142 844
<< m3 >>
rect 1098 800 1142 844
<< via2 >>
rect 1105 807 1135 837
<< m2 >>
rect 1479 800 1523 844
<< m3 >>
rect 1479 800 1523 844
<< via2 >>
rect 1486 807 1516 837
<< m2 >>
rect 1479 798 1523 842
<< m3 >>
rect 1479 798 1523 842
<< via2 >>
rect 1486 805 1516 835
<< m3 >>
rect 1106 925 1308 955
<< m2 >>
rect 1106 924 1136 955
<< m3 >>
rect 1103 924 1136 954
<< m2 >>
rect 1103 805 1133 954
<< m3 >>
rect 1101 805 1133 835
<< m2 >>
rect 1101 820 1131 835
<< m2 >>
rect 1099 918 1143 962
<< m3 >>
rect 1099 918 1143 962
<< via2 >>
rect 1106 925 1136 955
<< m2 >>
rect 1099 917 1143 961
<< m3 >>
rect 1099 917 1143 961
<< via2 >>
rect 1106 924 1136 954
<< m2 >>
rect 1096 917 1140 961
<< m3 >>
rect 1096 917 1140 961
<< via2 >>
rect 1103 924 1133 954
<< m2 >>
rect 1096 798 1140 842
<< m3 >>
rect 1096 798 1140 842
<< via2 >>
rect 1103 805 1133 835
<< m2 >>
rect 1094 813 1138 842
<< m3 >>
rect 1094 813 1138 842
<< via2 >>
rect 1101 820 1131 835
<< m2 >>
rect 1101 1220 1131 1235
<< m2 >>
rect 1101 805 1131 1235
<< m2 >>
rect 1101 805 1131 820
<< m2 >>
rect 1677 1220 1707 1235
<< m2 >>
rect 1677 808 1707 1235
<< m2 >>
rect 1677 808 1707 838
<< m2 >>
rect 1677 406 1707 838
<< m2 >>
rect 1677 406 1707 436
<< m2 >>
rect 1677 405 1707 436
<< m2 >>
rect 1677 405 1707 435
<< m2 >>
rect 1677 420 1707 435
<< m3 >>
rect 1104 1085 1500 1115
<< m2 >>
rect 1104 803 1134 1115
<< m3 >>
rect 1101 803 1134 833
<< m2 >>
rect 1101 420 1131 833
<< m2 >>
rect 1097 1078 1141 1122
<< m3 >>
rect 1097 1078 1141 1122
<< via2 >>
rect 1104 1085 1134 1115
<< m2 >>
rect 1097 796 1141 840
<< m3 >>
rect 1097 796 1141 840
<< via2 >>
rect 1104 803 1134 833
<< m2 >>
rect 1094 796 1138 840
<< m3 >>
rect 1094 796 1138 840
<< via2 >>
rect 1101 803 1131 833
<< m2 >>
rect 1485 1084 1515 1100
<< m3 >>
rect 1108 1084 1515 1114
<< m2 >>
rect 1108 926 1138 1114
<< m3 >>
rect 1107 926 1138 956
<< m2 >>
rect 1107 812 1137 956
<< m3 >>
rect 1106 812 1137 842
<< m2 >>
rect 1106 807 1136 842
<< m3 >>
rect 1101 807 1136 837
<< m2 >>
rect 1101 805 1131 837
<< m3 >>
rect 1116 805 1131 835
<< m2 >>
rect 1478 1077 1522 1107
<< m3 >>
rect 1478 1077 1522 1107
<< via2 >>
rect 1485 1084 1515 1100
<< m2 >>
rect 1101 1077 1145 1121
<< m3 >>
rect 1101 1077 1145 1121
<< via2 >>
rect 1108 1084 1138 1114
<< m2 >>
rect 1101 919 1145 963
<< m3 >>
rect 1101 919 1145 963
<< via2 >>
rect 1108 926 1138 956
<< m2 >>
rect 1100 919 1144 963
<< m3 >>
rect 1100 919 1144 963
<< via2 >>
rect 1107 926 1137 956
<< m2 >>
rect 1100 805 1144 849
<< m3 >>
rect 1100 805 1144 849
<< via2 >>
rect 1107 812 1137 842
<< m2 >>
rect 1099 805 1143 849
<< m3 >>
rect 1099 805 1143 849
<< via2 >>
rect 1106 812 1136 842
<< m2 >>
rect 1099 800 1143 844
<< m3 >>
rect 1099 800 1143 844
<< via2 >>
rect 1106 807 1136 837
<< m2 >>
rect 1094 800 1138 844
<< m3 >>
rect 1094 800 1138 844
<< via2 >>
rect 1101 807 1131 837
<< m2 >>
rect 1109 798 1138 842
<< m3 >>
rect 1109 798 1138 842
<< via2 >>
rect 1116 805 1131 835
<< m3 >>
rect 1293 285 1500 315
<< m2 >>
rect 1293 140 1323 315
<< m2 >>
rect 1286 278 1330 322
<< m3 >>
rect 1286 278 1330 322
<< via2 >>
rect 1293 285 1323 315
<< m2 >>
rect 1485 300 1515 316
<< m3 >>
rect 1101 286 1515 316
<< m2 >>
rect 1101 286 1131 420
<< m2 >>
rect 1478 293 1522 323
<< m3 >>
rect 1478 293 1522 323
<< via2 >>
rect 1485 300 1515 316
<< m2 >>
rect 1094 279 1138 323
<< m3 >>
rect 1094 279 1138 323
<< via2 >>
rect 1101 286 1131 316
<< m2 >>
rect 1485 300 1515 315
<< m3 >>
rect 1295 285 1515 315
<< m2 >>
rect 1295 285 1325 1556
<< m3 >>
rect 1293 1526 1325 1556
<< m2 >>
rect 1293 1526 1323 2140
<< m2 >>
rect 1478 293 1522 322
<< m3 >>
rect 1478 293 1522 322
<< via2 >>
rect 1485 300 1515 315
<< m2 >>
rect 1288 278 1332 322
<< m3 >>
rect 1288 278 1332 322
<< via2 >>
rect 1295 285 1325 315
<< m2 >>
rect 1288 1519 1332 1563
<< m3 >>
rect 1288 1519 1332 1563
<< via2 >>
rect 1295 1526 1325 1556
<< m2 >>
rect 1286 1519 1330 1563
<< m3 >>
rect 1286 1519 1330 1563
<< via2 >>
rect 1293 1526 1323 1556
<< m2 >>
rect 1485 300 1515 834
<< m2 >>
rect 1485 804 1515 834
<< m2 >>
rect 1485 804 1515 1236
<< m2 >>
rect 1485 1206 1515 1236
<< m2 >>
rect 1485 1206 1515 1836
<< m2 >>
rect 1485 1806 1515 1836
<< m2 >>
rect 1485 1806 1515 2300
<< m2 >>
rect 1485 300 1515 315
<< m2 >>
rect 1485 285 1515 715
<< m2 >>
rect 1485 685 1515 700
<< m2 >>
rect 1485 300 1515 433
<< m2 >>
rect 1485 403 1515 433
<< m2 >>
rect 1485 403 1515 713
<< m2 >>
rect 1485 683 1515 713
<< m2 >>
rect 1485 683 1515 700
<< m2 >>
rect 1485 300 1515 315
<< m3 >>
rect 1107 285 1515 315
<< m2 >>
rect 1107 285 1137 831
<< m3 >>
rect 1101 801 1137 831
<< m2 >>
rect 1101 801 1131 820
<< m2 >>
rect 1478 293 1522 322
<< m3 >>
rect 1478 293 1522 322
<< via2 >>
rect 1485 300 1515 315
<< m2 >>
rect 1100 278 1144 322
<< m3 >>
rect 1100 278 1144 322
<< via2 >>
rect 1107 285 1137 315
<< m2 >>
rect 1100 794 1144 838
<< m3 >>
rect 1100 794 1144 838
<< via2 >>
rect 1107 801 1137 831
<< m2 >>
rect 1094 794 1138 827
<< m3 >>
rect 1094 794 1138 827
<< via2 >>
rect 1101 801 1131 820
<< m2 >>
rect 1293 140 1323 312
<< m3 >>
rect 1293 282 1324 312
<< m2 >>
rect 1294 282 1324 551
<< m3 >>
rect 1294 521 1326 551
<< m2 >>
rect 1296 521 1326 713
<< m3 >>
rect 1296 683 1512 713
<< m2 >>
rect 1482 683 1512 714
<< m3 >>
rect 1482 684 1514 714
<< m2 >>
rect 1484 684 1514 715
<< m3 >>
rect 1484 685 1500 715
<< m2 >>
rect 1286 275 1330 319
<< m3 >>
rect 1286 275 1330 319
<< via2 >>
rect 1293 282 1323 312
<< m2 >>
rect 1287 275 1331 319
<< m3 >>
rect 1287 275 1331 319
<< via2 >>
rect 1294 282 1324 312
<< m2 >>
rect 1287 514 1331 558
<< m3 >>
rect 1287 514 1331 558
<< via2 >>
rect 1294 521 1324 551
<< m2 >>
rect 1289 514 1333 558
<< m3 >>
rect 1289 514 1333 558
<< via2 >>
rect 1296 521 1326 551
<< m2 >>
rect 1289 676 1333 720
<< m3 >>
rect 1289 676 1333 720
<< via2 >>
rect 1296 683 1326 713
<< m2 >>
rect 1475 676 1519 720
<< m3 >>
rect 1475 676 1519 720
<< via2 >>
rect 1482 683 1512 713
<< m2 >>
rect 1475 677 1519 721
<< m3 >>
rect 1475 677 1519 721
<< via2 >>
rect 1482 684 1512 714
<< m2 >>
rect 1477 677 1521 721
<< m3 >>
rect 1477 677 1521 721
<< via2 >>
rect 1484 684 1514 714
<< m2 >>
rect 1477 678 1507 722
<< m3 >>
rect 1477 678 1507 722
<< via2 >>
rect 1484 685 1500 715
<< m2 >>
rect 1101 420 1131 710
<< m3 >>
rect 1101 680 1511 710
<< m2 >>
rect 1481 680 1511 713
<< m3 >>
rect 1481 683 1515 713
<< m2 >>
rect 1485 683 1515 700
<< m2 >>
rect 1094 673 1138 717
<< m3 >>
rect 1094 673 1138 717
<< via2 >>
rect 1101 680 1131 710
<< m2 >>
rect 1474 673 1518 717
<< m3 >>
rect 1474 673 1518 717
<< via2 >>
rect 1481 680 1511 710
<< m2 >>
rect 1474 676 1518 720
<< m3 >>
rect 1474 676 1518 720
<< via2 >>
rect 1481 683 1511 713
<< m2 >>
rect 1478 676 1522 707
<< m3 >>
rect 1478 676 1522 707
<< via2 >>
rect 1485 683 1515 700
<< m2 >>
rect 1005 300 1035 709
<< m3 >>
rect 1005 679 1036 709
<< m2 >>
rect 1006 679 1036 828
<< m3 >>
rect 1006 798 1127 828
<< m2 >>
rect 1097 798 1127 832
<< m3 >>
rect 1097 802 1131 832
<< m2 >>
rect 1101 802 1131 820
<< m2 >>
rect 998 672 1042 716
<< m3 >>
rect 998 672 1042 716
<< via2 >>
rect 1005 679 1035 709
<< m2 >>
rect 999 672 1043 716
<< m3 >>
rect 999 672 1043 716
<< via2 >>
rect 1006 679 1036 709
<< m2 >>
rect 999 791 1043 835
<< m3 >>
rect 999 791 1043 835
<< via2 >>
rect 1006 798 1036 828
<< m2 >>
rect 1090 791 1134 835
<< m3 >>
rect 1090 791 1134 835
<< via2 >>
rect 1097 798 1127 828
<< m2 >>
rect 1090 795 1134 839
<< m3 >>
rect 1090 795 1134 839
<< via2 >>
rect 1097 802 1127 832
<< m2 >>
rect 1094 795 1138 827
<< m3 >>
rect 1094 795 1138 827
<< via2 >>
rect 1101 802 1131 820
<< m2 >>
rect 1101 2526 1131 2820
<< m3 >>
rect 1101 2526 1611 2556
<< m2 >>
rect 1581 2525 1611 2556
<< m3 >>
rect 1581 2525 1884 2555
<< m2 >>
rect 1094 2519 1138 2563
<< m3 >>
rect 1094 2519 1138 2563
<< via2 >>
rect 1101 2526 1131 2556
<< m2 >>
rect 1574 2519 1618 2563
<< m3 >>
rect 1574 2519 1618 2563
<< via2 >>
rect 1581 2526 1611 2556
<< m2 >>
rect 1574 2518 1618 2562
<< m3 >>
rect 1574 2518 1618 2562
<< via2 >>
rect 1581 2525 1611 2555
<< m3 >>
rect 1116 2805 1513 2835
<< m2 >>
rect 1483 2805 1513 2835
<< m3 >>
rect 1483 2805 1515 2835
<< m2 >>
rect 1485 2805 1515 2835
<< m3 >>
rect 1485 2805 1692 2835
<< m2 >>
rect 1476 2798 1520 2842
<< m3 >>
rect 1476 2798 1520 2842
<< via2 >>
rect 1483 2805 1513 2835
<< m2 >>
rect 1476 2798 1520 2842
<< m3 >>
rect 1476 2798 1520 2842
<< via2 >>
rect 1483 2805 1513 2835
<< m2 >>
rect 1478 2798 1522 2842
<< m3 >>
rect 1478 2798 1522 2842
<< via2 >>
rect 1485 2805 1515 2835
<< m2 >>
rect 1478 2798 1522 2842
<< m3 >>
rect 1478 2798 1522 2842
<< via2 >>
rect 1485 2805 1515 2835
<< m2 >>
rect 1101 2820 1131 2835
<< m2 >>
rect 1101 2405 1131 2835
<< m2 >>
rect 1101 2405 1131 2420
<< m2 >>
rect 1101 2804 1131 2820
<< m3 >>
rect 1101 2804 1133 2834
<< m2 >>
rect 1103 2405 1133 2834
<< m3 >>
rect 1103 2405 1515 2435
<< m2 >>
rect 1485 2405 1515 2435
<< m3 >>
rect 1485 2405 1692 2435
<< m2 >>
rect 1094 2797 1138 2827
<< m3 >>
rect 1094 2797 1138 2827
<< via2 >>
rect 1101 2804 1131 2820
<< m2 >>
rect 1096 2797 1140 2841
<< m3 >>
rect 1096 2797 1140 2841
<< via2 >>
rect 1103 2804 1133 2834
<< m2 >>
rect 1096 2398 1140 2442
<< m3 >>
rect 1096 2398 1140 2442
<< via2 >>
rect 1103 2405 1133 2435
<< m2 >>
rect 1478 2398 1522 2442
<< m3 >>
rect 1478 2398 1522 2442
<< via2 >>
rect 1485 2405 1515 2435
<< m2 >>
rect 1478 2398 1522 2442
<< m3 >>
rect 1478 2398 1522 2442
<< via2 >>
rect 1485 2405 1515 2435
<< m3 >>
rect 1106 2685 1500 2715
<< m2 >>
rect 1106 2525 1136 2715
<< m3 >>
rect 1105 2525 1136 2555
<< m2 >>
rect 1105 2407 1135 2555
<< m3 >>
rect 1102 2407 1135 2437
<< m2 >>
rect 1102 2405 1132 2437
<< m3 >>
rect 1116 2405 1132 2435
<< m2 >>
rect 1099 2678 1143 2722
<< m3 >>
rect 1099 2678 1143 2722
<< via2 >>
rect 1106 2685 1136 2715
<< m2 >>
rect 1099 2518 1143 2562
<< m3 >>
rect 1099 2518 1143 2562
<< via2 >>
rect 1106 2525 1136 2555
<< m2 >>
rect 1098 2518 1142 2562
<< m3 >>
rect 1098 2518 1142 2562
<< via2 >>
rect 1105 2525 1135 2555
<< m2 >>
rect 1098 2400 1142 2444
<< m3 >>
rect 1098 2400 1142 2444
<< via2 >>
rect 1105 2407 1135 2437
<< m2 >>
rect 1095 2400 1139 2444
<< m3 >>
rect 1095 2400 1139 2444
<< via2 >>
rect 1102 2407 1132 2437
<< m2 >>
rect 1109 2398 1139 2442
<< m3 >>
rect 1109 2398 1139 2442
<< via2 >>
rect 1116 2405 1132 2435
<< m2 >>
rect 1677 2420 1707 2820
<< m2 >>
rect 1293 2140 1323 2433
<< m3 >>
rect 1293 2403 1706 2433
<< m2 >>
rect 1676 2403 1706 2435
<< m3 >>
rect 1676 2405 1692 2435
<< m2 >>
rect 1286 2396 1330 2440
<< m3 >>
rect 1286 2396 1330 2440
<< via2 >>
rect 1293 2403 1323 2433
<< m2 >>
rect 1669 2396 1713 2440
<< m3 >>
rect 1669 2396 1713 2440
<< via2 >>
rect 1676 2403 1706 2433
<< m2 >>
rect 1669 2398 1699 2442
<< m3 >>
rect 1669 2398 1699 2442
<< via2 >>
rect 1676 2405 1692 2435
<< m2 >>
rect 1101 2420 1131 2435
<< m3 >>
rect 1101 2405 1321 2435
<< m2 >>
rect 1291 2405 1321 2435
<< m3 >>
rect 1291 2405 1707 2435
<< m2 >>
rect 1677 2405 1707 2420
<< m2 >>
rect 1094 2413 1138 2442
<< m3 >>
rect 1094 2413 1138 2442
<< via2 >>
rect 1101 2420 1131 2435
<< m2 >>
rect 1284 2398 1328 2442
<< m3 >>
rect 1284 2398 1328 2442
<< via2 >>
rect 1291 2405 1321 2435
<< m2 >>
rect 1284 2398 1328 2442
<< m3 >>
rect 1284 2398 1328 2442
<< via2 >>
rect 1291 2405 1321 2435
<< m2 >>
rect 1670 2398 1714 2427
<< m3 >>
rect 1670 2398 1714 2427
<< via2 >>
rect 1677 2405 1707 2420
<< labels >>
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 VSS
port 1 nsew signal bidirectional
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 VDD
port 2 nsew signal bidirectional
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 VIP
port 3 nsew signal bidirectional
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 VIN
port 4 nsew signal bidirectional
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 VO
port 5 nsew signal bidirectional
flabel  s 0 0 0 0 0 FreeSans 400 0 0 0 I_BIAS
port 6 nsew signal bidirectional
<< properties >>
<< end >>
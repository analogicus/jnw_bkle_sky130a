magic
tech sky130A
magscale 1 1
timestamp 1746013120
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4010
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWTR_CAPX1 None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 9048 0 1 500
box 0 0 540 540
use JNWATR_PCH_4C5F0 None_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7496 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 7496 0 1 4010
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 8072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP4<1>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 8072 0 1 4650
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 14250
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN1<5>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 14650
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT mirror1_MN1<5>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 14010
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN1<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4250
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 2072 0 1 4650
box 0 0 576 240
use JNWTR_RPPO8 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2300
box 0 0 1372 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 940 1720
use AALMISC_PNP_W3p40L3p40 load1_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2742 0 1 3180
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<0> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2072 0 1 3180
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<1> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2072 0 1 1170
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<2> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2742 0 1 1170
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<3> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2072 0 1 1840
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<4> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2742 0 1 1840
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<5> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2742 0 1 2510
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<6> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2072 0 1 2510
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<7> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 2072 0 1 500
box 0 0 670 670
<< locali >>
rect 100 15000 9788 15050
<< locali >>
rect 100 100 9788 150
<< m1 >>
rect 100 150 150 15000
<< m1 >>
rect 9738 150 9788 15000
<< locali >>
rect 93 14993 157 15057
<< m1 >>
rect 93 14993 157 15057
<< viali >>
rect 100 15000 150 15050
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 9731 14993 9795 15057
<< m1 >>
rect 9731 14993 9795 15057
<< viali >>
rect 9738 15000 9788 15050
<< locali >>
rect 9731 93 9795 157
<< m1 >>
rect 9731 93 9795 157
<< viali >>
rect 9738 100 9788 150
<< locali >>
rect 0 15100 9888 15150
<< locali >>
rect 0 0 9888 50
<< m1 >>
rect 0 50 50 15100
<< m1 >>
rect 9838 50 9888 15100
<< locali >>
rect -7 15093 57 15157
<< m1 >>
rect -7 15093 57 15157
<< viali >>
rect 0 15100 50 15150
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 9831 15093 9895 15157
<< m1 >>
rect 9831 15093 9895 15157
<< viali >>
rect 9838 15100 9888 15150
<< locali >>
rect 9831 -7 9895 57
<< m1 >>
rect 9831 -7 9895 57
<< viali >>
rect 9838 0 9888 50
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 7448 4550 7736 4590
<< locali >>
rect 7832 4430 7992 4470
<< locali >>
rect 8024 4550 8312 4590
<< locali >>
rect 8408 4430 8568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 14550 2312 14590
<< locali >>
rect 2408 14430 2568 14470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< locali >>
rect 2408 4430 2568 4470
<< locali >>
rect 2024 4550 2312 4590
<< m1 >>
rect 1872 100 1922 15050
<< m1 >>
rect 16046 100 16096 15050
<< locali >>
rect 1872 4082 16096 4178
<< locali >>
rect 16039 93 16103 157
<< m1 >>
rect 16039 93 16103 157
<< viali >>
rect 16046 100 16096 150
<< locali >>
rect 16039 14993 16103 15057
<< m1 >>
rect 16039 14993 16103 15057
<< viali >>
rect 16046 15000 16096 15050
<< locali >>
rect 1865 93 1929 157
<< m1 >>
rect 1865 93 1929 157
<< viali >>
rect 1872 100 1922 150
<< locali >>
rect 1865 14993 1929 15057
<< m1 >>
rect 1865 14993 1929 15057
<< viali >>
rect 1872 15000 1922 15050
<< locali >>
rect 1865 4075 1929 4185
<< m1 >>
rect 1865 4075 1929 4185
<< viali >>
rect 1872 4082 1922 4178
<< locali >>
rect 16039 4075 16103 4185
<< m1 >>
rect 16039 4075 16103 4185
<< viali >>
rect 16046 4082 16096 4178
<< locali >>
rect 16039 4075 16103 4185
<< m1 >>
rect 16039 4075 16103 4185
<< viali >>
rect 16046 4082 16096 4178
<< m1 >>
rect 1772 0 1822 15150
<< m1 >>
rect 2898 0 2948 15150
<< locali >>
rect 1772 14722 2948 14818
<< locali >>
rect 2891 -7 2955 57
<< m1 >>
rect 2891 -7 2955 57
<< viali >>
rect 2898 0 2948 50
<< locali >>
rect 2891 15093 2955 15157
<< m1 >>
rect 2891 15093 2955 15157
<< viali >>
rect 2898 15100 2948 15150
<< locali >>
rect 1765 -7 1829 57
<< m1 >>
rect 1765 -7 1829 57
<< viali >>
rect 1772 0 1822 50
<< locali >>
rect 1765 15093 1829 15157
<< m1 >>
rect 1765 15093 1829 15157
<< viali >>
rect 1772 15100 1822 15150
<< locali >>
rect 1765 14715 1829 14825
<< m1 >>
rect 1765 14715 1829 14825
<< viali >>
rect 1772 14722 1822 14818
<< locali >>
rect 2891 14715 2955 14825
<< m1 >>
rect 2891 14715 2955 14825
<< viali >>
rect 2898 14722 2948 14818
<< locali >>
rect 2891 14715 2955 14825
<< m1 >>
rect 2891 14715 2955 14825
<< viali >>
rect 2898 14722 2948 14818
<< m1 >>
rect 1772 0 1822 15150
<< m1 >>
rect 2898 0 2948 15150
<< locali >>
rect 1772 14082 2948 14178
<< locali >>
rect 2891 -7 2955 57
<< m1 >>
rect 2891 -7 2955 57
<< viali >>
rect 2898 0 2948 50
<< locali >>
rect 2891 15093 2955 15157
<< m1 >>
rect 2891 15093 2955 15157
<< viali >>
rect 2898 15100 2948 15150
<< locali >>
rect 1765 -7 1829 57
<< m1 >>
rect 1765 -7 1829 57
<< viali >>
rect 1772 0 1822 50
<< locali >>
rect 1765 15093 1829 15157
<< m1 >>
rect 1765 15093 1829 15157
<< viali >>
rect 1772 15100 1822 15150
<< locali >>
rect 1765 14075 1829 14185
<< m1 >>
rect 1765 14075 1829 14185
<< viali >>
rect 1772 14082 1822 14178
<< locali >>
rect 2891 14075 2955 14185
<< m1 >>
rect 2891 14075 2955 14185
<< viali >>
rect 2898 14082 2948 14178
<< locali >>
rect 2891 14075 2955 14185
<< m1 >>
rect 2891 14075 2955 14185
<< viali >>
rect 2898 14082 2948 14178
<< locali >>
rect 0 3964 1372 4020
<< locali >>
rect -7 3957 57 4027
<< m1 >>
rect -7 3957 57 4027
<< viali >>
rect 0 3964 50 4020
<< locali >>
rect 1315 3957 1379 4027
<< m1 >>
rect 1315 3957 1379 4027
<< viali >>
rect 1322 3964 1372 4020
<< locali >>
rect 0 2300 1372 2356
<< locali >>
rect -7 2293 57 2363
<< m1 >>
rect -7 2293 57 2363
<< viali >>
rect 0 2300 50 2356
<< locali >>
rect 1315 2293 1379 2363
<< m1 >>
rect 1315 2293 1379 2363
<< viali >>
rect 1322 2300 1372 2356
<< locali >>
rect 0 2164 940 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 883 2157 947 2227
<< m1 >>
rect 883 2157 947 2227
<< viali >>
rect 890 2164 940 2220
<< locali >>
rect 0 500 940 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 883 493 947 563
<< m1 >>
rect 883 493 947 563
<< viali >>
rect 890 500 940 556
use OTA U1_OTA 
transform 1 0 9938 0 1 0
box 0 0 4438 6440
<< labels >>
flabel locali s 100 15000 9788 15050 0 FreeSans 400 0 0 0 VDD
port 4 nsew signal bidirectional
flabel locali s 0 15100 9888 15150 0 FreeSans 400 0 0 0 VSS
port 5 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1745837706
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5740
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWTR_CAPX1 None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4740
box 0 0 540 540
use JNWATR_PCH_4C5F0 None_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5980
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6380
box 0 0 576 240
use JNWTR_RPPO8 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2320
box 0 0 1372 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 600 0 1 500
box 0 0 940 1720
use AALMISC_PNP_W3p40L3p40 load1_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 1154 0 1 8150
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<0> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 12260
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<1> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 1154 0 1 12260
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<2> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 1154 0 1 10890
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<3> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 10890
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<4> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 1154 0 1 9520
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<5> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 1154 0 1 6780
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<6> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6780
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<7> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 8150
box 0 0 670 670
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< m3 >>
rect 629 5993 739 6047
<< via2 >>
rect 636 6000 732 6040
<< via1 >>
rect 636 6000 732 6040
<< locali >>
rect 775 1953 933 2087
<< m1 >>
rect 775 1953 933 2087
<< m2 >>
rect 775 1953 933 2087
<< m3 >>
rect 775 1953 933 2087
<< via2 >>
rect 782 1960 926 2080
<< via1 >>
rect 782 1960 926 2080
<< viali >>
rect 782 1960 926 2080
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< m3 >>
rect 373 6153 419 6207
<< via2 >>
rect 380 6160 412 6200
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< locali >>
rect 1424 8456 1562 8522
<< m1 >>
rect 1424 8456 1562 8522
<< m2 >>
rect 1424 8456 1562 8522
<< m3 >>
rect 1424 8456 1562 8522
<< via2 >>
rect 1431 8463 1555 8515
<< via1 >>
rect 1431 8463 1555 8515
<< viali >>
rect 1431 8463 1555 8515
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< m2 >>
rect 475 3773 633 3907
<< m3 >>
rect 475 3773 633 3907
<< via2 >>
rect 482 3780 626 3900
<< via1 >>
rect 482 3780 626 3900
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 1207 1953 1365 2087
<< m1 >>
rect 1207 1953 1365 2087
<< m2 >>
rect 1207 1953 1365 2087
<< m3 >>
rect 1207 1953 1365 2087
<< via2 >>
rect 1214 1960 1358 2080
<< via1 >>
rect 1214 1960 1358 2080
<< viali >>
rect 1214 1960 1358 2080
<< m3 >>
rect 663 5795 693 6018
<< m2 >>
rect 663 5795 869 5825
<< m3 >>
rect 839 4867 869 5825
<< m2 >>
rect 839 4867 1013 4897
<< m3 >>
rect 983 2595 1013 4897
<< m2 >>
rect 839 2595 1013 2625
<< m3 >>
rect 839 2018 869 2625
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< locali >>
rect 775 1953 933 2087
<< m1 >>
rect 775 1953 933 2087
<< viali >>
rect 782 1960 926 2080
<< m2 >>
rect 656 5788 700 5832
<< m3 >>
rect 656 5788 700 5832
<< via2 >>
rect 663 5795 693 5825
<< m2 >>
rect 832 5788 876 5832
<< m3 >>
rect 832 5788 876 5832
<< via2 >>
rect 839 5795 869 5825
<< m2 >>
rect 832 4860 876 4904
<< m3 >>
rect 832 4860 876 4904
<< via2 >>
rect 839 4867 869 4897
<< m2 >>
rect 976 4860 1020 4904
<< m3 >>
rect 976 4860 1020 4904
<< via2 >>
rect 983 4867 1013 4897
<< m2 >>
rect 976 2588 1020 2632
<< m3 >>
rect 976 2588 1020 2632
<< via2 >>
rect 983 2595 1013 2625
<< m2 >>
rect 832 2588 876 2632
<< m3 >>
rect 832 2588 876 2632
<< via2 >>
rect 839 2595 869 2625
<< m3 >>
rect 375 4963 405 6178
<< m2 >>
rect 375 4963 581 4993
<< m3 >>
rect 551 4754 581 4993
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m1 >>
rect 373 6153 419 6207
<< m2 >>
rect 373 6153 419 6207
<< via1 >>
rect 380 6160 412 6200
<< m2 >>
rect 368 4956 412 5000
<< m3 >>
rect 368 4956 412 5000
<< via2 >>
rect 375 4963 405 4993
<< m2 >>
rect 544 4956 588 5000
<< m3 >>
rect 544 4956 588 5000
<< via2 >>
rect 551 4963 581 4993
<< m2 >>
rect 678 6003 885 6033
<< m3 >>
rect 855 6003 885 6449
<< m2 >>
rect 855 6419 1045 6449
<< m3 >>
rect 1015 6419 1045 6593
<< m2 >>
rect 1015 6563 1189 6593
<< m3 >>
rect 1159 6563 1189 6737
<< m2 >>
rect 1159 6707 1333 6737
<< m3 >>
rect 1303 6707 1333 8129
<< m2 >>
rect 1303 8099 1509 8129
<< m3 >>
rect 1479 8099 1509 8482
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< m1 >>
rect 629 5993 739 6047
<< m2 >>
rect 629 5993 739 6047
<< via1 >>
rect 636 6000 732 6040
<< locali >>
rect 1424 8456 1562 8522
<< m1 >>
rect 1424 8456 1562 8522
<< viali >>
rect 1431 8463 1555 8515
<< m2 >>
rect 848 5996 892 6040
<< m3 >>
rect 848 5996 892 6040
<< via2 >>
rect 855 6003 885 6033
<< m2 >>
rect 848 6412 892 6456
<< m3 >>
rect 848 6412 892 6456
<< via2 >>
rect 855 6419 885 6449
<< m2 >>
rect 1008 6412 1052 6456
<< m3 >>
rect 1008 6412 1052 6456
<< via2 >>
rect 1015 6419 1045 6449
<< m2 >>
rect 1008 6556 1052 6600
<< m3 >>
rect 1008 6556 1052 6600
<< via2 >>
rect 1015 6563 1045 6593
<< m2 >>
rect 1152 6556 1196 6600
<< m3 >>
rect 1152 6556 1196 6600
<< via2 >>
rect 1159 6563 1189 6593
<< m2 >>
rect 1152 6700 1196 6744
<< m3 >>
rect 1152 6700 1196 6744
<< via2 >>
rect 1159 6707 1189 6737
<< m2 >>
rect 1296 6700 1340 6744
<< m3 >>
rect 1296 6700 1340 6744
<< via2 >>
rect 1303 6707 1333 6737
<< m2 >>
rect 1296 8092 1340 8136
<< m3 >>
rect 1296 8092 1340 8136
<< via2 >>
rect 1303 8099 1333 8129
<< m2 >>
rect 1472 8092 1516 8136
<< m3 >>
rect 1472 8092 1516 8136
<< via2 >>
rect 1479 8099 1509 8129
<< m3 >>
rect 534 3569 564 3840
<< m2 >>
rect 534 3569 708 3599
<< m3 >>
rect 678 3409 708 3599
<< m2 >>
rect 678 3409 868 3439
<< m3 >>
rect 838 2849 868 3439
<< m2 >>
rect 838 2849 1124 2879
<< m3 >>
rect 1094 2257 1124 2879
<< m2 >>
rect 1094 2257 1300 2287
<< m3 >>
rect 1270 2016 1300 2287
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 1207 1953 1365 2087
<< m1 >>
rect 1207 1953 1365 2087
<< viali >>
rect 1214 1960 1358 2080
<< m2 >>
rect 527 3562 571 3606
<< m3 >>
rect 527 3562 571 3606
<< via2 >>
rect 534 3569 564 3599
<< m2 >>
rect 671 3562 715 3606
<< m3 >>
rect 671 3562 715 3606
<< via2 >>
rect 678 3569 708 3599
<< m2 >>
rect 671 3402 715 3446
<< m3 >>
rect 671 3402 715 3446
<< via2 >>
rect 678 3409 708 3439
<< m2 >>
rect 831 3402 875 3446
<< m3 >>
rect 831 3402 875 3446
<< via2 >>
rect 838 3409 868 3439
<< m2 >>
rect 831 2842 875 2886
<< m3 >>
rect 831 2842 875 2886
<< via2 >>
rect 838 2849 868 2879
<< m2 >>
rect 1087 2842 1131 2886
<< m3 >>
rect 1087 2842 1131 2886
<< via2 >>
rect 1094 2849 1124 2879
<< m2 >>
rect 1087 2250 1131 2294
<< m3 >>
rect 1087 2250 1131 2294
<< via2 >>
rect 1094 2257 1124 2287
<< m2 >>
rect 1263 2250 1307 2294
<< m3 >>
rect 1263 2250 1307 2294
<< via2 >>
rect 1270 2257 1300 2287
<< locali >>
rect 100 13280 2024 13330
<< locali >>
rect 100 100 2024 150
<< m1 >>
rect 100 150 150 13280
<< m1 >>
rect 1974 150 2024 13280
<< locali >>
rect 93 13273 157 13337
<< m1 >>
rect 93 13273 157 13337
<< viali >>
rect 100 13280 150 13330
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1967 13273 2031 13337
<< m1 >>
rect 1967 13273 2031 13337
<< viali >>
rect 1974 13280 2024 13330
<< locali >>
rect 1967 93 2031 157
<< m1 >>
rect 1967 93 2031 157
<< viali >>
rect 1974 100 2024 150
<< locali >>
rect 0 13380 2124 13430
<< locali >>
rect 0 0 2124 50
<< m1 >>
rect 0 50 50 13380
<< m1 >>
rect 2074 50 2124 13380
<< locali >>
rect -7 13373 57 13437
<< m1 >>
rect -7 13373 57 13437
<< viali >>
rect 0 13380 50 13430
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2067 13373 2131 13437
<< m1 >>
rect 2067 13373 2131 13437
<< viali >>
rect 2074 13380 2124 13430
<< locali >>
rect 2067 -7 2131 57
<< m1 >>
rect 2067 -7 2131 57
<< viali >>
rect 2074 0 2124 50
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 636 6160 796 6200
<< locali >>
rect 252 6280 540 6320
<< locali >>
rect 100 5812 2024 5908
<< locali >>
rect 93 5805 157 5915
<< m1 >>
rect 93 5805 157 5915
<< viali >>
rect 100 5812 150 5908
<< locali >>
rect 1967 5805 2031 5915
<< m1 >>
rect 1967 5805 2031 5915
<< viali >>
rect 1974 5812 2024 5908
<< locali >>
rect 0 3984 2124 4040
<< locali >>
rect -7 3977 57 4047
<< m1 >>
rect -7 3977 57 4047
<< viali >>
rect 0 3984 50 4040
<< locali >>
rect 2067 3977 2131 4047
<< m1 >>
rect 2067 3977 2131 4047
<< viali >>
rect 2074 3984 2124 4040
<< locali >>
rect 0 2320 2124 2376
<< locali >>
rect -7 2313 57 2383
<< m1 >>
rect -7 2313 57 2383
<< viali >>
rect 0 2320 50 2376
<< locali >>
rect 2067 2313 2131 2383
<< m1 >>
rect 2067 2313 2131 2383
<< viali >>
rect 2074 2320 2124 2376
<< locali >>
rect 0 2164 2124 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 2067 2157 2131 2227
<< m1 >>
rect 2067 2157 2131 2227
<< viali >>
rect 2074 2164 2124 2220
<< locali >>
rect 0 500 2124 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 2067 493 2131 563
<< m1 >>
rect 2067 493 2131 563
<< viali >>
rect 2074 500 2124 556
use OTA U1_OTA 
transform 1 0 2174 0 1 21970
box 0 0 5322 8490
<< labels >>
flabel locali s 100 13280 2024 13330 0 FreeSans 400 0 0 0 VDD
port 31 nsew signal bidirectional
flabel locali s 0 13380 2124 13430 0 FreeSans 400 0 0 0 VSS
port 32 nsew signal bidirectional
flabel m1 s 636 6000 732 6040 0 FreeSans 400 0 0 0 OUT
port 33 nsew signal bidirectional
<< properties >>
<< end >>
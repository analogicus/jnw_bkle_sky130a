magic
tech sky130A
magscale 1 1
timestamp 1744203138
<< checkpaint >>
rect 0 0 0 0
use COMP2 U1_COMP2 
transform 1 0 4500 0 1 0
box -450 -650 1602 3850
use OTA_Manuel U2_OTA_Manuel 
transform 1 0 6552 0 1 0
box -600 -800 3820 4400
<< labels >>
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1748586004
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0  diff1_MP3<3> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 504
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  diff1_MP3<3>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 264
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP3<2> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  diff1_MP3<2>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP3<1> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 1304
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<0> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 1304
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<3> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  diff1_MP4<3>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 2504
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP4<2> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 2104
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  diff1_MP4<2>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 2504
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP4<1> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<0> ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 1704
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror1_MP2 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 904
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror1_MP1 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 904
box 0 0 576 400
use JNWATR_NCH_4C5F0  mirror2_MN1 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 3304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 3704
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 868 0 1 3064
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN2 ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 3304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 3704
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748586004
transform 1 0 292 0 1 3064
box 0 0 576 240
use JNWTR_RPPO16  bias1_RH1 ../JNW_TR_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 4104
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH2 ../JNW_TR_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 5874
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH3 ../JNW_TR_SKY130A
timestamp 1748586004
transform 1 0 200 0 1 7644
box 0 0 2236 1720
<< m2 >>
rect 388 1486 979 1516
<< m2 >>
rect 821 1486 979 1516
<< m3 >>
rect 821 686 851 1516
<< m2 >>
rect 821 686 979 716
<< m2 >>
rect 388 686 979 716
<< m2 >>
rect 814 1479 858 1523
<< m3 >>
rect 814 1479 858 1523
<< via2 >>
rect 821 1486 851 1516
<< m2 >>
rect 814 679 858 723
<< m3 >>
rect 814 679 858 723
<< via2 >>
rect 821 686 851 716
<< m2 >>
rect 821 2286 964 2316
<< m3 >>
rect 821 1886 851 2316
<< m2 >>
rect 821 1886 979 1916
<< m2 >>
rect 373 1886 979 1916
<< m2 >>
rect 245 1886 403 1916
<< m3 >>
rect 245 1886 275 2316
<< m2 >>
rect 245 2286 388 2316
<< m2 >>
rect 814 2279 858 2323
<< m3 >>
rect 814 2279 858 2323
<< via2 >>
rect 821 2286 851 2316
<< m2 >>
rect 814 1879 858 1923
<< m3 >>
rect 814 1879 858 1923
<< via2 >>
rect 821 1886 851 1916
<< m2 >>
rect 238 1879 282 1923
<< m3 >>
rect 238 1879 282 1923
<< via2 >>
rect 245 1886 275 1916
<< m2 >>
rect 238 2279 282 2323
<< m3 >>
rect 238 2279 282 2323
<< via2 >>
rect 245 2286 275 2316
<< m3 >>
rect 661 2127 691 3342
<< m3 >>
rect 661 1727 691 2157
<< m2 >>
rect 661 1727 1267 1757
<< m3 >>
rect 1237 1727 1267 2142
<< m2 >>
rect 654 1720 698 1764
<< m3 >>
rect 654 1720 698 1764
<< via2 >>
rect 661 1727 691 1757
<< m2 >>
rect 1230 1720 1274 1764
<< m3 >>
rect 1230 1720 1274 1764
<< via2 >>
rect 1237 1727 1267 1757
<< m2 >>
rect 388 3487 979 3517
<< m2 >>
rect 949 3487 1411 3517
<< m3 >>
rect 1381 1327 1411 3517
<< m2 >>
rect 661 1327 1411 1357
<< m2 >>
rect 661 1327 1267 1357
<< m2 >>
rect 1237 1327 1411 1357
<< m3 >>
rect 1381 527 1411 1357
<< m2 >>
rect 1237 527 1411 557
<< m2 >>
rect 676 527 1267 557
<< m2 >>
rect 1374 3480 1418 3524
<< m3 >>
rect 1374 3480 1418 3524
<< via2 >>
rect 1381 3487 1411 3517
<< m2 >>
rect 1374 1320 1418 1364
<< m3 >>
rect 1374 1320 1418 1364
<< via2 >>
rect 1381 1327 1411 1357
<< m2 >>
rect 1374 1320 1418 1364
<< m3 >>
rect 1374 1320 1418 1364
<< via2 >>
rect 1381 1327 1411 1357
<< m2 >>
rect 1374 520 1418 564
<< m3 >>
rect 1374 520 1418 564
<< via2 >>
rect 1381 527 1411 557
<< m2 >>
rect 261 921 676 951
<< m3 >>
rect 261 921 291 1639
<< m2 >>
rect 261 1609 499 1639
<< m2 >>
rect 149 1609 499 1639
<< m3 >>
rect 149 1609 179 2039
<< m2 >>
rect 149 2009 499 2039
<< m2 >>
rect 149 2009 499 2039
<< m3 >>
rect 149 2009 179 2439
<< m2 >>
rect 149 2409 499 2439
<< m2 >>
rect 469 2409 1075 2439
<< m2 >>
rect 1045 2409 1507 2439
<< m3 >>
rect 1477 2009 1507 2439
<< m2 >>
rect 1045 2009 1507 2039
<< m2 >>
rect 1045 2009 1507 2039
<< m3 >>
rect 1477 1609 1507 2039
<< m2 >>
rect 1045 1609 1507 1639
<< m2 >>
rect 1045 1609 1507 1639
<< m3 >>
rect 1477 809 1507 1639
<< m2 >>
rect 1045 809 1507 839
<< m2 >>
rect 484 809 1075 839
<< m2 >>
rect 254 914 298 958
<< m3 >>
rect 254 914 298 958
<< via2 >>
rect 261 921 291 951
<< m2 >>
rect 254 1602 298 1646
<< m3 >>
rect 254 1602 298 1646
<< via2 >>
rect 261 1609 291 1639
<< m2 >>
rect 142 1602 186 1646
<< m3 >>
rect 142 1602 186 1646
<< via2 >>
rect 149 1609 179 1639
<< m2 >>
rect 142 2002 186 2046
<< m3 >>
rect 142 2002 186 2046
<< via2 >>
rect 149 2009 179 2039
<< m2 >>
rect 142 2002 186 2046
<< m3 >>
rect 142 2002 186 2046
<< via2 >>
rect 149 2009 179 2039
<< m2 >>
rect 142 2402 186 2446
<< m3 >>
rect 142 2402 186 2446
<< via2 >>
rect 149 2409 179 2439
<< m2 >>
rect 1470 2402 1514 2446
<< m3 >>
rect 1470 2402 1514 2446
<< via2 >>
rect 1477 2409 1507 2439
<< m2 >>
rect 1470 2002 1514 2046
<< m3 >>
rect 1470 2002 1514 2046
<< via2 >>
rect 1477 2009 1507 2039
<< m2 >>
rect 1470 2002 1514 2046
<< m3 >>
rect 1470 2002 1514 2046
<< via2 >>
rect 1477 2009 1507 2039
<< m2 >>
rect 1470 1602 1514 1646
<< m3 >>
rect 1470 1602 1514 1646
<< via2 >>
rect 1477 1609 1507 1639
<< m2 >>
rect 1470 1602 1514 1646
<< m3 >>
rect 1470 1602 1514 1646
<< via2 >>
rect 1477 1609 1507 1639
<< m2 >>
rect 1470 802 1514 846
<< m3 >>
rect 1470 802 1514 846
<< via2 >>
rect 1477 809 1507 839
<< m3 >>
rect 2165 1085 2195 5628
<< m2 >>
rect 949 1085 2195 1115
<< m2 >>
rect 388 1085 979 1115
<< m2 >>
rect 2158 1078 2202 1122
<< m3 >>
rect 2158 1078 2202 1122
<< via2 >>
rect 2165 1085 2195 1115
<< m3 >>
rect 438 5622 468 6869
<< m2 >>
rect 438 6839 2196 6869
<< m3 >>
rect 2166 6839 2196 7382
<< m2 >>
rect 431 6832 475 6876
<< m3 >>
rect 431 6832 475 6876
<< via2 >>
rect 438 6839 468 6869
<< m2 >>
rect 2159 6832 2203 6876
<< m3 >>
rect 2159 6832 2203 6876
<< via2 >>
rect 2166 6839 2196 6869
<< m3 >>
rect 438 7387 468 8938
<< m2 >>
rect 438 8908 2196 8938
<< m3 >>
rect 2166 8908 2196 9163
<< m2 >>
rect 431 8901 475 8945
<< m3 >>
rect 431 8901 475 8945
<< via2 >>
rect 438 8908 468 8938
<< m2 >>
rect 2159 8901 2203 8945
<< m3 >>
rect 2159 8901 2203 8945
<< via2 >>
rect 2166 8908 2196 8938
<< locali >>
rect 100 9414 2536 9464
<< locali >>
rect 100 100 2536 150
<< m1 >>
rect 100 150 150 9414
<< m1 >>
rect 2486 150 2536 9414
<< locali >>
rect 93 9407 157 9471
<< m1 >>
rect 93 9407 157 9471
<< viali >>
rect 100 9414 150 9464
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2479 9407 2543 9471
<< m1 >>
rect 2479 9407 2543 9471
<< viali >>
rect 2486 9414 2536 9464
<< locali >>
rect 2479 93 2543 157
<< m1 >>
rect 2479 93 2543 157
<< viali >>
rect 2486 100 2536 150
<< locali >>
rect 0 9514 2636 9564
<< locali >>
rect 0 0 2636 50
<< m1 >>
rect 0 50 50 9514
<< m1 >>
rect 2586 50 2636 9514
<< locali >>
rect -7 9507 57 9571
<< m1 >>
rect -7 9507 57 9571
<< viali >>
rect 0 9514 50 9564
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2579 9507 2643 9571
<< m1 >>
rect 2579 9507 2643 9571
<< viali >>
rect 2586 9514 2636 9564
<< locali >>
rect 2579 -7 2643 57
<< m1 >>
rect 2579 -7 2643 57
<< viali >>
rect 2586 0 2636 50
<< locali >>
rect 208 9104 526 9224
<< locali >>
rect 100 5768 2536 5824
<< locali >>
rect 93 5761 157 5831
<< m1 >>
rect 93 5761 157 5831
<< viali >>
rect 100 5768 150 5824
<< locali >>
rect 2479 5761 2543 5831
<< m1 >>
rect 2479 5761 2543 5831
<< viali >>
rect 2486 5768 2536 5824
<< locali >>
rect 100 4104 2536 4160
<< locali >>
rect 93 4097 157 4167
<< m1 >>
rect 93 4097 157 4167
<< viali >>
rect 100 4104 150 4160
<< locali >>
rect 2479 4097 2543 4167
<< m1 >>
rect 2479 4097 2543 4167
<< viali >>
rect 2486 4104 2536 4160
<< locali >>
rect 100 7538 2536 7594
<< locali >>
rect 93 7531 157 7601
<< m1 >>
rect 93 7531 157 7601
<< viali >>
rect 100 7538 150 7594
<< locali >>
rect 2479 7531 2543 7601
<< m1 >>
rect 2479 7531 2543 7601
<< viali >>
rect 2486 7538 2536 7594
<< locali >>
rect 100 5874 2536 5930
<< locali >>
rect 93 5867 157 5937
<< m1 >>
rect 93 5867 157 5937
<< viali >>
rect 100 5874 150 5930
<< locali >>
rect 2479 5867 2543 5937
<< m1 >>
rect 2479 5867 2543 5937
<< viali >>
rect 2486 5874 2536 5930
<< locali >>
rect 100 9308 2536 9364
<< locali >>
rect 93 9301 157 9371
<< m1 >>
rect 93 9301 157 9371
<< viali >>
rect 100 9308 150 9364
<< locali >>
rect 2479 9301 2543 9371
<< m1 >>
rect 2479 9301 2543 9371
<< viali >>
rect 2486 9308 2536 9364
<< locali >>
rect 100 7644 2536 7700
<< locali >>
rect 93 7637 157 7707
<< m1 >>
rect 93 7637 157 7707
<< viali >>
rect 100 7644 150 7700
<< locali >>
rect 2479 7637 2543 7707
<< m1 >>
rect 2479 7637 2543 7707
<< viali >>
rect 2486 7644 2536 7700
<< locali >>
rect 244 1204 532 1244
<< locali >>
rect 820 1204 1108 1244
<< locali >>
rect 1204 1084 1364 1124
<< locali >>
rect 820 3604 1108 3644
<< locali >>
rect 1204 3484 1364 3524
<< locali >>
rect 244 3604 532 3644
<< locali >>
rect 0 336 2636 432
<< locali >>
rect -7 329 57 439
<< m1 >>
rect -7 329 57 439
<< viali >>
rect 0 336 50 432
<< locali >>
rect 2579 329 2643 439
<< m1 >>
rect 2579 329 2643 439
<< viali >>
rect 2586 336 2636 432
<< locali >>
rect 0 2576 2636 2672
<< locali >>
rect -7 2569 57 2679
<< m1 >>
rect -7 2569 57 2679
<< viali >>
rect 0 2576 50 2672
<< locali >>
rect 2579 2569 2643 2679
<< m1 >>
rect 2579 2569 2643 2679
<< viali >>
rect 2586 2576 2636 2672
<< locali >>
rect 100 3776 2536 3872
<< locali >>
rect 93 3769 157 3879
<< m1 >>
rect 93 3769 157 3879
<< viali >>
rect 100 3776 150 3872
<< locali >>
rect 2479 3769 2543 3879
<< m1 >>
rect 2479 3769 2543 3879
<< viali >>
rect 2486 3776 2536 3872
<< locali >>
rect 100 3136 2536 3232
<< locali >>
rect 93 3129 157 3239
<< m1 >>
rect 93 3129 157 3239
<< viali >>
rect 100 3136 150 3232
<< locali >>
rect 2479 3129 2543 3239
<< m1 >>
rect 2479 3129 2543 3239
<< viali >>
rect 2486 3136 2536 3232
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 365 1477 411 1531
<< m2 >>
rect 365 1477 411 1531
<< via1 >>
rect 372 1484 404 1524
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 365 2277 411 2331
<< m2 >>
rect 365 2277 411 2331
<< via1 >>
rect 372 2284 404 2324
<< m1 >>
rect 941 2277 987 2331
<< m2 >>
rect 941 2277 987 2331
<< via1 >>
rect 948 2284 980 2324
<< m1 >>
rect 941 1877 987 1931
<< m2 >>
rect 941 1877 987 1931
<< via1 >>
rect 948 1884 980 1924
<< m1 >>
rect 941 1877 987 1931
<< m2 >>
rect 941 1877 987 1931
<< via1 >>
rect 948 1884 980 1924
<< m1 >>
rect 365 1877 411 1931
<< m2 >>
rect 365 1877 411 1931
<< via1 >>
rect 372 1884 404 1924
<< m1 >>
rect 365 1877 411 1931
<< m2 >>
rect 365 1877 411 1931
<< via1 >>
rect 372 1884 404 1924
<< m1 >>
rect 621 2117 731 2171
<< m2 >>
rect 621 2117 731 2171
<< m3 >>
rect 621 2117 731 2171
<< via2 >>
rect 628 2124 724 2164
<< via1 >>
rect 628 2124 724 2164
<< m1 >>
rect 621 2117 731 2171
<< m2 >>
rect 621 2117 731 2171
<< m3 >>
rect 621 2117 731 2171
<< via2 >>
rect 628 2124 724 2164
<< via1 >>
rect 628 2124 724 2164
<< m1 >>
rect 1197 2117 1307 2171
<< m2 >>
rect 1197 2117 1307 2171
<< m3 >>
rect 1197 2117 1307 2171
<< via2 >>
rect 1204 2124 1300 2164
<< via1 >>
rect 1204 2124 1300 2164
<< m1 >>
rect 1197 1717 1307 1771
<< m2 >>
rect 1197 1717 1307 1771
<< via1 >>
rect 1204 1724 1300 1764
<< m1 >>
rect 1197 1717 1307 1771
<< m2 >>
rect 1197 1717 1307 1771
<< m3 >>
rect 1197 1717 1307 1771
<< via2 >>
rect 1204 1724 1300 1764
<< via1 >>
rect 1204 1724 1300 1764
<< m1 >>
rect 621 1717 731 1771
<< m2 >>
rect 621 1717 731 1771
<< m3 >>
rect 621 1717 731 1771
<< via2 >>
rect 628 1724 724 1764
<< via1 >>
rect 628 1724 724 1764
<< m1 >>
rect 621 1717 731 1771
<< m2 >>
rect 621 1717 731 1771
<< via1 >>
rect 628 1724 724 1764
<< m1 >>
rect 621 3317 731 3371
<< m2 >>
rect 621 3317 731 3371
<< m3 >>
rect 621 3317 731 3371
<< via2 >>
rect 628 3324 724 3364
<< via1 >>
rect 628 3324 724 3364
<< m1 >>
rect 621 517 731 571
<< m2 >>
rect 621 517 731 571
<< via1 >>
rect 628 524 724 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 1197 517 1307 571
<< m2 >>
rect 1197 517 1307 571
<< via1 >>
rect 1204 524 1300 564
<< m1 >>
rect 621 1317 731 1371
<< m2 >>
rect 621 1317 731 1371
<< via1 >>
rect 628 1324 724 1364
<< m1 >>
rect 621 1317 731 1371
<< m2 >>
rect 621 1317 731 1371
<< via1 >>
rect 628 1324 724 1364
<< m1 >>
rect 1197 1317 1307 1371
<< m2 >>
rect 1197 1317 1307 1371
<< via1 >>
rect 1204 1324 1300 1364
<< m1 >>
rect 1197 1317 1307 1371
<< m2 >>
rect 1197 1317 1307 1371
<< via1 >>
rect 1204 1324 1300 1364
<< m1 >>
rect 1197 1317 1307 1371
<< m2 >>
rect 1197 1317 1307 1371
<< via1 >>
rect 1204 1324 1300 1364
<< m1 >>
rect 941 3477 987 3531
<< m2 >>
rect 941 3477 987 3531
<< via1 >>
rect 948 3484 980 3524
<< m1 >>
rect 941 3477 987 3531
<< m2 >>
rect 941 3477 987 3531
<< via1 >>
rect 948 3484 980 3524
<< m1 >>
rect 365 3477 411 3531
<< m2 >>
rect 365 3477 411 3531
<< via1 >>
rect 372 3484 404 3524
<< m1 >>
rect 429 797 539 851
<< m2 >>
rect 429 797 539 851
<< via1 >>
rect 436 804 532 844
<< m1 >>
rect 1005 797 1115 851
<< m2 >>
rect 1005 797 1115 851
<< via1 >>
rect 1012 804 1108 844
<< m1 >>
rect 1005 797 1115 851
<< m2 >>
rect 1005 797 1115 851
<< via1 >>
rect 1012 804 1108 844
<< m1 >>
rect 429 1597 539 1651
<< m2 >>
rect 429 1597 539 1651
<< via1 >>
rect 436 1604 532 1644
<< m1 >>
rect 429 1597 539 1651
<< m2 >>
rect 429 1597 539 1651
<< via1 >>
rect 436 1604 532 1644
<< m1 >>
rect 1005 1597 1115 1651
<< m2 >>
rect 1005 1597 1115 1651
<< via1 >>
rect 1012 1604 1108 1644
<< m1 >>
rect 1005 1597 1115 1651
<< m2 >>
rect 1005 1597 1115 1651
<< via1 >>
rect 1012 1604 1108 1644
<< m1 >>
rect 429 2397 539 2451
<< m2 >>
rect 429 2397 539 2451
<< via1 >>
rect 436 2404 532 2444
<< m1 >>
rect 429 2397 539 2451
<< m2 >>
rect 429 2397 539 2451
<< via1 >>
rect 436 2404 532 2444
<< m1 >>
rect 1005 2397 1115 2451
<< m2 >>
rect 1005 2397 1115 2451
<< via1 >>
rect 1012 2404 1108 2444
<< m1 >>
rect 1005 2397 1115 2451
<< m2 >>
rect 1005 2397 1115 2451
<< via1 >>
rect 1012 2404 1108 2444
<< m1 >>
rect 1005 1997 1115 2051
<< m2 >>
rect 1005 1997 1115 2051
<< via1 >>
rect 1012 2004 1108 2044
<< m1 >>
rect 1005 1997 1115 2051
<< m2 >>
rect 1005 1997 1115 2051
<< via1 >>
rect 1012 2004 1108 2044
<< m1 >>
rect 429 1997 539 2051
<< m2 >>
rect 429 1997 539 2051
<< via1 >>
rect 436 2004 532 2044
<< m1 >>
rect 429 1997 539 2051
<< m2 >>
rect 429 1997 539 2051
<< via1 >>
rect 436 2004 532 2044
<< m1 >>
rect 621 917 731 971
<< m2 >>
rect 621 917 731 971
<< via1 >>
rect 628 924 724 964
<< m1 >>
rect 365 1077 411 1131
<< m2 >>
rect 365 1077 411 1131
<< via1 >>
rect 372 1084 404 1124
<< m1 >>
rect 941 1077 987 1131
<< m2 >>
rect 941 1077 987 1131
<< via1 >>
rect 948 1084 980 1124
<< m1 >>
rect 941 1077 987 1131
<< m2 >>
rect 941 1077 987 1131
<< via1 >>
rect 948 1084 980 1124
<< locali >>
rect 2103 5557 2261 5691
<< m1 >>
rect 2103 5557 2261 5691
<< m2 >>
rect 2103 5557 2261 5691
<< m3 >>
rect 2103 5557 2261 5691
<< via2 >>
rect 2110 5564 2254 5684
<< via1 >>
rect 2110 5564 2254 5684
<< viali >>
rect 2110 5564 2254 5684
<< locali >>
rect 375 5557 533 5691
<< m1 >>
rect 375 5557 533 5691
<< m2 >>
rect 375 5557 533 5691
<< m3 >>
rect 375 5557 533 5691
<< via2 >>
rect 382 5564 526 5684
<< via1 >>
rect 382 5564 526 5684
<< viali >>
rect 382 5564 526 5684
<< locali >>
rect 2103 7327 2261 7461
<< m1 >>
rect 2103 7327 2261 7461
<< m2 >>
rect 2103 7327 2261 7461
<< m3 >>
rect 2103 7327 2261 7461
<< via2 >>
rect 2110 7334 2254 7454
<< via1 >>
rect 2110 7334 2254 7454
<< viali >>
rect 2110 7334 2254 7454
<< locali >>
rect 375 7327 533 7461
<< m1 >>
rect 375 7327 533 7461
<< m2 >>
rect 375 7327 533 7461
<< m3 >>
rect 375 7327 533 7461
<< via2 >>
rect 382 7334 526 7454
<< via1 >>
rect 382 7334 526 7454
<< viali >>
rect 382 7334 526 7454
<< locali >>
rect 2103 9097 2261 9231
<< m1 >>
rect 2103 9097 2261 9231
<< m2 >>
rect 2103 9097 2261 9231
<< m3 >>
rect 2103 9097 2261 9231
<< via2 >>
rect 2110 9104 2254 9224
<< via1 >>
rect 2110 9104 2254 9224
<< viali >>
rect 2110 9104 2254 9224
<< labels >>
flabel m2 s 388 1486 979 1516 0 FreeSans 400 0 0 0 IN+
port 74 nsew signal bidirectional
flabel m2 s 821 2286 964 2316 0 FreeSans 400 0 0 0 IN-
port 75 nsew signal bidirectional
flabel locali s 0 9514 2636 9564 0 FreeSans 400 0 0 0 VDD
port 76 nsew signal bidirectional
flabel locali s 100 9414 2536 9464 0 FreeSans 400 0 0 0 VSS
port 77 nsew signal bidirectional
flabel m3 s 661 2127 691 3342 0 FreeSans 400 0 0 0 OUT
port 78 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
timestamp 1729602094
<< metal3 >>
rect 0 0 340 340
<< mimcap >>
rect 20 310 320 320
rect 20 30 30 310
rect 310 30 320 310
rect 20 20 320 30
<< mimcapcontact >>
rect 30 30 310 310
<< metal4 >>
rect 0 310 340 340
rect 0 30 30 310
rect 310 30 340 310
rect 0 0 340 30
<< labels >>
flabel metal4 s 0 0 340 50 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel metal3 s 0 0 340 50 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 340 340
<< end >>

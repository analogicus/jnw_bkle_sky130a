magic
tech sky130A
magscale 1 1
timestamp 1746459945
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1800
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1800
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<1>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<0>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2600
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2600
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 3400
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 3400
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 -40
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 -40
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 3446
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 6986
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 5216
box 0 0 2236 1720
<< m1 >>
rect 941 1973 987 2027
<< m2 >>
rect 941 1973 987 2027
<< via1 >>
rect 948 1980 980 2020
<< m1 >>
rect 365 1973 411 2027
<< m2 >>
rect 365 1973 411 2027
<< via1 >>
rect 372 1980 404 2020
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< m3 >>
rect 365 1573 411 1627
<< via2 >>
rect 372 1580 404 1620
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< m3 >>
rect 941 1573 987 1627
<< via2 >>
rect 948 1580 980 1620
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< m3 >>
rect 365 2773 411 2827
<< via2 >>
rect 372 2780 404 2820
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< via1 >>
rect 948 2780 980 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< m3 >>
rect 941 2773 987 2827
<< via2 >>
rect 948 2780 980 2820
<< via1 >>
rect 948 2780 980 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< via1 >>
rect 948 2780 980 2820
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< m3 >>
rect 621 2213 731 2267
<< via2 >>
rect 628 2220 724 2260
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< m3 >>
rect 621 2213 731 2267
<< via2 >>
rect 628 2220 724 2260
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 1197 2213 1307 2267
<< m2 >>
rect 1197 2213 1307 2267
<< m3 >>
rect 1197 2213 1307 2267
<< via2 >>
rect 1204 2220 1300 2260
<< via1 >>
rect 1204 2220 1300 2260
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< m3 >>
rect 621 2613 731 2667
<< via2 >>
rect 628 2620 724 2660
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< m3 >>
rect 621 2613 731 2667
<< via2 >>
rect 628 2620 724 2660
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< m3 >>
rect 1197 2613 1307 2667
<< via2 >>
rect 1204 2620 1300 2660
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< m3 >>
rect 1197 2613 1307 2667
<< via2 >>
rect 1204 2620 1300 2660
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< m3 >>
rect 1197 1813 1307 1867
<< via2 >>
rect 1204 1820 1300 1860
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< m3 >>
rect 1197 1813 1307 1867
<< via2 >>
rect 1204 1820 1300 1860
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< m3 >>
rect 621 1813 731 1867
<< via2 >>
rect 628 1820 724 1860
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< m3 >>
rect 621 1813 731 1867
<< via2 >>
rect 628 1820 724 1860
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1413 731 1467
<< m2 >>
rect 621 1413 731 1467
<< m3 >>
rect 621 1413 731 1467
<< via2 >>
rect 628 1420 724 1460
<< via1 >>
rect 628 1420 724 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< m3 >>
rect 941 373 987 427
<< via2 >>
rect 948 380 980 420
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< m3 >>
rect 941 373 987 427
<< via2 >>
rect 948 380 980 420
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< m3 >>
rect 1197 213 1307 267
<< via2 >>
rect 1204 220 1300 260
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< m3 >>
rect 1197 213 1307 267
<< via2 >>
rect 1204 220 1300 260
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 365 373 411 427
<< m2 >>
rect 365 373 411 427
<< via1 >>
rect 372 380 404 420
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< m3 >>
rect 1005 2093 1115 2147
<< via2 >>
rect 1012 2100 1108 2140
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 429 2093 539 2147
<< m2 >>
rect 429 2093 539 2147
<< via1 >>
rect 436 2100 532 2140
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< m3 >>
rect 429 1693 539 1747
<< via2 >>
rect 436 1700 532 1740
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< m3 >>
rect 1005 1693 1115 1747
<< via2 >>
rect 1012 1700 1108 1740
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 429 2493 539 2547
<< m2 >>
rect 429 2493 539 2547
<< via1 >>
rect 436 2500 532 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< m3 >>
rect 1005 2493 1115 2547
<< via2 >>
rect 1012 2500 1108 2540
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 429 2893 539 2947
<< m2 >>
rect 429 2893 539 2947
<< m3 >>
rect 429 2893 539 2947
<< via2 >>
rect 436 2900 532 2940
<< via1 >>
rect 436 2900 532 2940
<< m1 >>
rect 429 2893 539 2947
<< m2 >>
rect 429 2893 539 2947
<< via1 >>
rect 436 2900 532 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< m3 >>
rect 1005 2893 1115 2947
<< via2 >>
rect 1012 2900 1108 2940
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 621 3013 731 3067
<< m2 >>
rect 621 3013 731 3067
<< via1 >>
rect 628 3020 724 3060
<< m1 >>
rect 365 3173 411 3227
<< m2 >>
rect 365 3173 411 3227
<< via1 >>
rect 372 3180 404 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< m3 >>
rect 941 3173 987 3227
<< via2 >>
rect 948 3180 980 3220
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< m3 >>
rect 941 3173 987 3227
<< via2 >>
rect 948 3180 980 3220
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< via1 >>
rect 1204 3020 1300 3060
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< m3 >>
rect 1197 3013 1307 3067
<< via2 >>
rect 1204 3020 1300 3060
<< via1 >>
rect 1204 3020 1300 3060
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< via1 >>
rect 1204 3020 1300 3060
<< locali >>
rect 2103 4899 2261 5033
<< m1 >>
rect 2103 4899 2261 5033
<< m2 >>
rect 2103 4899 2261 5033
<< m3 >>
rect 2103 4899 2261 5033
<< via2 >>
rect 2110 4906 2254 5026
<< via1 >>
rect 2110 4906 2254 5026
<< viali >>
rect 2110 4906 2254 5026
<< locali >>
rect 375 4899 533 5033
<< m1 >>
rect 375 4899 533 5033
<< m2 >>
rect 375 4899 533 5033
<< via1 >>
rect 382 4906 526 5026
<< viali >>
rect 382 4906 526 5026
<< locali >>
rect 2103 8439 2261 8573
<< m1 >>
rect 2103 8439 2261 8573
<< m2 >>
rect 2103 8439 2261 8573
<< via1 >>
rect 2110 8446 2254 8566
<< viali >>
rect 2110 8446 2254 8566
<< locali >>
rect 375 8439 533 8573
<< m1 >>
rect 375 8439 533 8573
<< m2 >>
rect 375 8439 533 8573
<< via1 >>
rect 382 8446 526 8566
<< viali >>
rect 382 8446 526 8566
<< locali >>
rect 2103 6669 2261 6803
<< m1 >>
rect 2103 6669 2261 6803
<< m2 >>
rect 2103 6669 2261 6803
<< via1 >>
rect 2110 6676 2254 6796
<< viali >>
rect 2110 6676 2254 6796
<< m2 >>
rect 243 1982 386 2012
<< m3 >>
rect 243 1582 273 2012
<< m2 >>
rect 243 1582 401 1612
<< m3 >>
rect 371 1582 401 1612
<< m2 >>
rect 371 1582 977 1612
<< m3 >>
rect 947 1582 977 1612
<< m2 >>
rect 819 1582 977 1612
<< m3 >>
rect 819 1582 849 2012
<< m2 >>
rect 819 1982 962 2012
<< m1 >>
rect 941 1973 987 2027
<< m2 >>
rect 941 1973 987 2027
<< via1 >>
rect 948 1980 980 2020
<< m1 >>
rect 365 1973 411 2027
<< m2 >>
rect 365 1973 411 2027
<< via1 >>
rect 372 1980 404 2020
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m2 >>
rect 236 1975 280 2019
<< m3 >>
rect 236 1975 280 2019
<< via2 >>
rect 243 1982 273 2012
<< m2 >>
rect 236 1575 280 1619
<< m3 >>
rect 236 1575 280 1619
<< via2 >>
rect 243 1582 273 1612
<< m2 >>
rect 364 1575 408 1619
<< m3 >>
rect 364 1575 408 1619
<< via2 >>
rect 371 1582 401 1612
<< m2 >>
rect 364 1575 408 1619
<< m3 >>
rect 364 1575 408 1619
<< via2 >>
rect 371 1582 401 1612
<< m2 >>
rect 940 1575 984 1619
<< m3 >>
rect 940 1575 984 1619
<< via2 >>
rect 947 1582 977 1612
<< m2 >>
rect 940 1575 984 1619
<< m3 >>
rect 940 1575 984 1619
<< via2 >>
rect 947 1582 977 1612
<< m2 >>
rect 812 1575 856 1619
<< m3 >>
rect 812 1575 856 1619
<< via2 >>
rect 819 1582 849 1612
<< m2 >>
rect 812 1975 856 2019
<< m3 >>
rect 812 1975 856 2019
<< via2 >>
rect 819 1982 849 2012
<< m2 >>
rect 819 2382 962 2412
<< m3 >>
rect 819 2382 849 2812
<< m2 >>
rect 819 2782 977 2812
<< m3 >>
rect 947 2782 977 2812
<< m2 >>
rect 371 2782 977 2812
<< m3 >>
rect 371 2782 401 2812
<< m2 >>
rect 243 2782 401 2812
<< m3 >>
rect 243 2382 273 2812
<< m2 >>
rect 243 2382 386 2412
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 365 2773 411 2827
<< m2 >>
rect 365 2773 411 2827
<< via1 >>
rect 372 2780 404 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< via1 >>
rect 948 2780 980 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< via1 >>
rect 948 2780 980 2820
<< m1 >>
rect 941 2773 987 2827
<< m2 >>
rect 941 2773 987 2827
<< via1 >>
rect 948 2780 980 2820
<< m2 >>
rect 812 2375 856 2419
<< m3 >>
rect 812 2375 856 2419
<< via2 >>
rect 819 2382 849 2412
<< m2 >>
rect 812 2775 856 2819
<< m3 >>
rect 812 2775 856 2819
<< via2 >>
rect 819 2782 849 2812
<< m2 >>
rect 940 2775 984 2819
<< m3 >>
rect 940 2775 984 2819
<< via2 >>
rect 947 2782 977 2812
<< m2 >>
rect 940 2775 984 2819
<< m3 >>
rect 940 2775 984 2819
<< via2 >>
rect 947 2782 977 2812
<< m2 >>
rect 364 2775 408 2819
<< m3 >>
rect 364 2775 408 2819
<< via2 >>
rect 371 2782 401 2812
<< m2 >>
rect 364 2775 408 2819
<< m3 >>
rect 364 2775 408 2819
<< via2 >>
rect 371 2782 401 2812
<< m2 >>
rect 236 2775 280 2819
<< m3 >>
rect 236 2775 280 2819
<< via2 >>
rect 243 2782 273 2812
<< m2 >>
rect 236 2375 280 2419
<< m3 >>
rect 236 2375 280 2419
<< via2 >>
rect 243 2382 273 2412
<< m2 >>
rect 147 223 674 253
<< m3 >>
rect 147 223 177 2253
<< m2 >>
rect 147 2223 689 2253
<< m3 >>
rect 659 2223 689 2253
<< m3 >>
rect 659 2223 689 2653
<< m3 >>
rect 659 2623 689 2653
<< m2 >>
rect 659 2623 1265 2653
<< m3 >>
rect 1235 2623 1265 2653
<< m3 >>
rect 1235 2238 1265 2653
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< via1 >>
rect 628 2220 724 2260
<< m1 >>
rect 1197 2213 1307 2267
<< m2 >>
rect 1197 2213 1307 2267
<< via1 >>
rect 1204 2220 1300 2260
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 621 2613 731 2667
<< m2 >>
rect 621 2613 731 2667
<< via1 >>
rect 628 2620 724 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 1197 2613 1307 2667
<< m2 >>
rect 1197 2613 1307 2667
<< via1 >>
rect 1204 2620 1300 2660
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< via1 >>
rect 628 220 724 260
<< m2 >>
rect 140 216 184 260
<< m3 >>
rect 140 216 184 260
<< via2 >>
rect 147 223 177 253
<< m2 >>
rect 140 2216 184 2260
<< m3 >>
rect 140 2216 184 2260
<< via2 >>
rect 147 2223 177 2253
<< m2 >>
rect 652 2216 696 2260
<< m3 >>
rect 652 2216 696 2260
<< via2 >>
rect 659 2223 689 2253
<< m2 >>
rect 652 2616 696 2660
<< m3 >>
rect 652 2616 696 2660
<< via2 >>
rect 659 2623 689 2653
<< m2 >>
rect 1228 2616 1272 2660
<< m3 >>
rect 1228 2616 1272 2660
<< via2 >>
rect 1235 2623 1265 2653
<< m2 >>
rect 387 383 978 413
<< m3 >>
rect 948 383 978 413
<< m3 >>
rect 948 223 978 413
<< m2 >>
rect 948 223 1266 253
<< m3 >>
rect 1236 223 1266 253
<< m3 >>
rect 1236 223 1266 1453
<< m3 >>
rect 1236 1423 1266 1453
<< m3 >>
rect 1236 1423 1266 1853
<< m3 >>
rect 1236 1823 1266 1853
<< m2 >>
rect 660 1823 1266 1853
<< m3 >>
rect 660 1823 690 1853
<< m3 >>
rect 660 1438 690 1853
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 1197 1813 1307 1867
<< m2 >>
rect 1197 1813 1307 1867
<< via1 >>
rect 1204 1820 1300 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1813 731 1867
<< m2 >>
rect 621 1813 731 1867
<< via1 >>
rect 628 1820 724 1860
<< m1 >>
rect 621 1413 731 1467
<< m2 >>
rect 621 1413 731 1467
<< via1 >>
rect 628 1420 724 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< via1 >>
rect 1204 220 1300 260
<< m1 >>
rect 365 373 411 427
<< m2 >>
rect 365 373 411 427
<< via1 >>
rect 372 380 404 420
<< m2 >>
rect 941 376 985 420
<< m3 >>
rect 941 376 985 420
<< via2 >>
rect 948 383 978 413
<< m2 >>
rect 941 216 985 260
<< m3 >>
rect 941 216 985 260
<< via2 >>
rect 948 223 978 253
<< m2 >>
rect 1229 216 1273 260
<< m3 >>
rect 1229 216 1273 260
<< via2 >>
rect 1236 223 1266 253
<< m2 >>
rect 1229 1816 1273 1860
<< m3 >>
rect 1229 1816 1273 1860
<< via2 >>
rect 1236 1823 1266 1853
<< m2 >>
rect 653 1816 697 1860
<< m3 >>
rect 653 1816 697 1860
<< via2 >>
rect 660 1823 690 1853
<< m2 >>
rect 500 3017 675 3047
<< m3 >>
rect 500 2633 530 3047
<< m2 >>
rect 340 2633 530 2663
<< m3 >>
rect 340 2505 370 2663
<< m2 >>
rect 340 2505 498 2535
<< m2 >>
rect 516 2905 1074 2935
<< m3 >>
rect 1044 2905 1074 2935
<< m2 >>
rect 1044 2905 1410 2935
<< m3 >>
rect 1380 2505 1410 2935
<< m2 >>
rect 1044 2505 1410 2535
<< m3 >>
rect 1044 2505 1074 2535
<< m2 >>
rect 1044 2505 1410 2535
<< m3 >>
rect 1380 2105 1410 2535
<< m2 >>
rect 1044 2105 1410 2135
<< m3 >>
rect 1044 2105 1074 2135
<< m2 >>
rect 1044 2105 1410 2135
<< m3 >>
rect 1380 1705 1410 2135
<< m2 >>
rect 1044 1705 1410 1735
<< m3 >>
rect 1044 1705 1074 1735
<< m2 >>
rect 468 1705 1074 1735
<< m3 >>
rect 468 1705 498 1735
<< m2 >>
rect 52 1705 498 1735
<< m3 >>
rect 52 1705 82 2135
<< m2 >>
rect 52 2105 483 2135
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 1005 2093 1115 2147
<< m2 >>
rect 1005 2093 1115 2147
<< via1 >>
rect 1012 2100 1108 2140
<< m1 >>
rect 429 2093 539 2147
<< m2 >>
rect 429 2093 539 2147
<< via1 >>
rect 436 2100 532 2140
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 429 1693 539 1747
<< m2 >>
rect 429 1693 539 1747
<< via1 >>
rect 436 1700 532 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 1005 1693 1115 1747
<< m2 >>
rect 1005 1693 1115 1747
<< via1 >>
rect 1012 1700 1108 1740
<< m1 >>
rect 429 2493 539 2547
<< m2 >>
rect 429 2493 539 2547
<< via1 >>
rect 436 2500 532 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 1005 2493 1115 2547
<< m2 >>
rect 1005 2493 1115 2547
<< via1 >>
rect 1012 2500 1108 2540
<< m1 >>
rect 429 2893 539 2947
<< m2 >>
rect 429 2893 539 2947
<< via1 >>
rect 436 2900 532 2940
<< m1 >>
rect 429 2893 539 2947
<< m2 >>
rect 429 2893 539 2947
<< via1 >>
rect 436 2900 532 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 1005 2893 1115 2947
<< m2 >>
rect 1005 2893 1115 2947
<< via1 >>
rect 1012 2900 1108 2940
<< m1 >>
rect 621 3013 731 3067
<< m2 >>
rect 621 3013 731 3067
<< via1 >>
rect 628 3020 724 3060
<< m2 >>
rect 493 3010 537 3054
<< m3 >>
rect 493 3010 537 3054
<< via2 >>
rect 500 3017 530 3047
<< m2 >>
rect 493 2626 537 2670
<< m3 >>
rect 493 2626 537 2670
<< via2 >>
rect 500 2633 530 2663
<< m2 >>
rect 333 2626 377 2670
<< m3 >>
rect 333 2626 377 2670
<< via2 >>
rect 340 2633 370 2663
<< m2 >>
rect 333 2498 377 2542
<< m3 >>
rect 333 2498 377 2542
<< via2 >>
rect 340 2505 370 2535
<< m2 >>
rect 1037 2898 1081 2942
<< m3 >>
rect 1037 2898 1081 2942
<< via2 >>
rect 1044 2905 1074 2935
<< m2 >>
rect 1037 2898 1081 2942
<< m3 >>
rect 1037 2898 1081 2942
<< via2 >>
rect 1044 2905 1074 2935
<< m2 >>
rect 1373 2898 1417 2942
<< m3 >>
rect 1373 2898 1417 2942
<< via2 >>
rect 1380 2905 1410 2935
<< m2 >>
rect 1373 2498 1417 2542
<< m3 >>
rect 1373 2498 1417 2542
<< via2 >>
rect 1380 2505 1410 2535
<< m2 >>
rect 1037 2498 1081 2542
<< m3 >>
rect 1037 2498 1081 2542
<< via2 >>
rect 1044 2505 1074 2535
<< m2 >>
rect 1037 2498 1081 2542
<< m3 >>
rect 1037 2498 1081 2542
<< via2 >>
rect 1044 2505 1074 2535
<< m2 >>
rect 1373 2498 1417 2542
<< m3 >>
rect 1373 2498 1417 2542
<< via2 >>
rect 1380 2505 1410 2535
<< m2 >>
rect 1373 2098 1417 2142
<< m3 >>
rect 1373 2098 1417 2142
<< via2 >>
rect 1380 2105 1410 2135
<< m2 >>
rect 1037 2098 1081 2142
<< m3 >>
rect 1037 2098 1081 2142
<< via2 >>
rect 1044 2105 1074 2135
<< m2 >>
rect 1037 2098 1081 2142
<< m3 >>
rect 1037 2098 1081 2142
<< via2 >>
rect 1044 2105 1074 2135
<< m2 >>
rect 1373 2098 1417 2142
<< m3 >>
rect 1373 2098 1417 2142
<< via2 >>
rect 1380 2105 1410 2135
<< m2 >>
rect 1373 1698 1417 1742
<< m3 >>
rect 1373 1698 1417 1742
<< via2 >>
rect 1380 1705 1410 1735
<< m2 >>
rect 1037 1698 1081 1742
<< m3 >>
rect 1037 1698 1081 1742
<< via2 >>
rect 1044 1705 1074 1735
<< m2 >>
rect 1037 1698 1081 1742
<< m3 >>
rect 1037 1698 1081 1742
<< via2 >>
rect 1044 1705 1074 1735
<< m2 >>
rect 461 1698 505 1742
<< m3 >>
rect 461 1698 505 1742
<< via2 >>
rect 468 1705 498 1735
<< m2 >>
rect 461 1698 505 1742
<< m3 >>
rect 461 1698 505 1742
<< via2 >>
rect 468 1705 498 1735
<< m2 >>
rect 45 1698 89 1742
<< m3 >>
rect 45 1698 89 1742
<< via2 >>
rect 52 1705 82 1735
<< m2 >>
rect 45 2098 89 2142
<< m3 >>
rect 45 2098 89 2142
<< via2 >>
rect 52 2105 82 2135
<< m3 >>
rect 2163 3019 2193 4970
<< m2 >>
rect 1235 3019 2193 3049
<< m3 >>
rect 1235 3019 1265 3049
<< m2 >>
rect 947 3019 1265 3049
<< m3 >>
rect 947 3019 977 3209
<< m3 >>
rect 947 3179 977 3209
<< m2 >>
rect 386 3179 977 3209
<< m1 >>
rect 365 3173 411 3227
<< m2 >>
rect 365 3173 411 3227
<< via1 >>
rect 372 3180 404 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 941 3173 987 3227
<< m2 >>
rect 941 3173 987 3227
<< via1 >>
rect 948 3180 980 3220
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< via1 >>
rect 1204 3020 1300 3060
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< via1 >>
rect 1204 3020 1300 3060
<< m1 >>
rect 1197 3013 1307 3067
<< m2 >>
rect 1197 3013 1307 3067
<< via1 >>
rect 1204 3020 1300 3060
<< locali >>
rect 2103 4899 2261 5033
<< m1 >>
rect 2103 4899 2261 5033
<< viali >>
rect 2110 4906 2254 5026
<< m2 >>
rect 2156 3012 2200 3056
<< m3 >>
rect 2156 3012 2200 3056
<< via2 >>
rect 2163 3019 2193 3049
<< m2 >>
rect 1228 3012 1272 3056
<< m3 >>
rect 1228 3012 1272 3056
<< via2 >>
rect 1235 3019 1265 3049
<< m2 >>
rect 1228 3012 1272 3056
<< m3 >>
rect 1228 3012 1272 3056
<< via2 >>
rect 1235 3019 1265 3049
<< m2 >>
rect 940 3012 984 3056
<< m3 >>
rect 940 3012 984 3056
<< via2 >>
rect 947 3019 977 3049
<< m2 >>
rect 940 3172 984 3216
<< m3 >>
rect 940 3172 984 3216
<< via2 >>
rect 947 3179 977 3209
<< m2 >>
rect 449 4950 2064 4980
<< m3 >>
rect 2034 4950 2064 8516
<< m2 >>
rect 2034 8486 2177 8516
<< locali >>
rect 375 4899 533 5033
<< m1 >>
rect 375 4899 533 5033
<< viali >>
rect 382 4906 526 5026
<< locali >>
rect 2103 8439 2261 8573
<< m1 >>
rect 2103 8439 2261 8573
<< viali >>
rect 2110 8446 2254 8566
<< m2 >>
rect 2027 4943 2071 4987
<< m3 >>
rect 2027 4943 2071 4987
<< via2 >>
rect 2034 4950 2064 4980
<< m2 >>
rect 2027 8479 2071 8523
<< m3 >>
rect 2027 8479 2071 8523
<< via2 >>
rect 2034 8486 2064 8516
<< m2 >>
rect 449 8488 1760 8518
<< m3 >>
rect 1730 6712 1760 8518
<< m2 >>
rect 1730 6712 2177 6742
<< locali >>
rect 375 8439 533 8573
<< m1 >>
rect 375 8439 533 8573
<< viali >>
rect 382 8446 526 8566
<< locali >>
rect 2103 6669 2261 6803
<< m1 >>
rect 2103 6669 2261 6803
<< viali >>
rect 2110 6676 2254 6796
<< m2 >>
rect 1723 8481 1767 8525
<< m3 >>
rect 1723 8481 1767 8525
<< via2 >>
rect 1730 8488 1760 8518
<< m2 >>
rect 1723 6705 1767 6749
<< m3 >>
rect 1723 6705 1767 6749
<< via2 >>
rect 1730 6712 1760 6742
<< locali >>
rect 100 8756 2536 8806
<< locali >>
rect 100 100 2536 150
<< m1 >>
rect 100 150 150 8756
<< m1 >>
rect 2486 150 2536 8756
<< locali >>
rect 93 8749 157 8813
<< m1 >>
rect 93 8749 157 8813
<< viali >>
rect 100 8756 150 8806
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2479 8749 2543 8813
<< m1 >>
rect 2479 8749 2543 8813
<< viali >>
rect 2486 8756 2536 8806
<< locali >>
rect 2479 93 2543 157
<< m1 >>
rect 2479 93 2543 157
<< viali >>
rect 2486 100 2536 150
<< locali >>
rect 0 8856 2636 8906
<< locali >>
rect 0 0 2636 50
<< m1 >>
rect 0 50 50 8856
<< m1 >>
rect 2586 50 2636 8856
<< locali >>
rect -7 8849 57 8913
<< m1 >>
rect -7 8849 57 8913
<< viali >>
rect 0 8856 50 8906
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2579 8849 2643 8913
<< m1 >>
rect 2579 8849 2643 8913
<< viali >>
rect 2586 8856 2636 8906
<< locali >>
rect 2579 -7 2643 57
<< m1 >>
rect 2579 -7 2643 57
<< viali >>
rect 2586 0 2636 50
<< locali >>
rect 208 6676 526 6796
<< locali >>
rect 100 5110 2536 5166
<< locali >>
rect 93 5103 157 5173
<< m1 >>
rect 93 5103 157 5173
<< viali >>
rect 100 5110 150 5166
<< locali >>
rect 2479 5103 2543 5173
<< m1 >>
rect 2479 5103 2543 5173
<< viali >>
rect 2486 5110 2536 5166
<< locali >>
rect 100 3446 2536 3502
<< locali >>
rect 93 3439 157 3509
<< m1 >>
rect 93 3439 157 3509
<< viali >>
rect 100 3446 150 3502
<< locali >>
rect 2479 3439 2543 3509
<< m1 >>
rect 2479 3439 2543 3509
<< viali >>
rect 2486 3446 2536 3502
<< locali >>
rect 100 8650 2536 8706
<< locali >>
rect 93 8643 157 8713
<< m1 >>
rect 93 8643 157 8713
<< viali >>
rect 100 8650 150 8706
<< locali >>
rect 2479 8643 2543 8713
<< m1 >>
rect 2479 8643 2543 8713
<< viali >>
rect 2486 8650 2536 8706
<< locali >>
rect 100 6986 2536 7042
<< locali >>
rect 93 6979 157 7049
<< m1 >>
rect 93 6979 157 7049
<< viali >>
rect 100 6986 150 7042
<< locali >>
rect 2479 6979 2543 7049
<< m1 >>
rect 2479 6979 2543 7049
<< viali >>
rect 2486 6986 2536 7042
<< locali >>
rect 100 6880 2536 6936
<< locali >>
rect 93 6873 157 6943
<< m1 >>
rect 93 6873 157 6943
<< viali >>
rect 100 6880 150 6936
<< locali >>
rect 2479 6873 2543 6943
<< m1 >>
rect 2479 6873 2543 6943
<< viali >>
rect 2486 6880 2536 6936
<< locali >>
rect 100 5216 2536 5272
<< locali >>
rect 93 5209 157 5279
<< m1 >>
rect 93 5209 157 5279
<< viali >>
rect 100 5216 150 5272
<< locali >>
rect 2479 5209 2543 5279
<< m1 >>
rect 2479 5209 2543 5279
<< viali >>
rect 2486 5216 2536 5272
<< locali >>
rect 244 3300 532 3340
<< locali >>
rect 820 3300 1108 3340
<< locali >>
rect 1204 3180 1364 3220
<< locali >>
rect 820 500 1108 540
<< locali >>
rect 1204 380 1364 420
<< locali >>
rect 244 500 532 540
<< locali >>
rect 0 1232 2636 1328
<< locali >>
rect -7 1225 57 1335
<< m1 >>
rect -7 1225 57 1335
<< viali >>
rect 0 1232 50 1328
<< locali >>
rect 2579 1225 2643 1335
<< m1 >>
rect 2579 1225 2643 1335
<< viali >>
rect 2586 1232 2636 1328
<< locali >>
rect 0 3472 2636 3568
<< locali >>
rect -7 3465 57 3575
<< m1 >>
rect -7 3465 57 3575
<< viali >>
rect 0 3472 50 3568
<< locali >>
rect 2579 3465 2643 3575
<< m1 >>
rect 2579 3465 2643 3575
<< viali >>
rect 2586 3472 2636 3568
<< locali >>
rect 100 672 2536 768
<< locali >>
rect 93 665 157 775
<< m1 >>
rect 93 665 157 775
<< viali >>
rect 100 672 150 768
<< locali >>
rect 2479 665 2543 775
<< m1 >>
rect 2479 665 2543 775
<< viali >>
rect 2486 672 2536 768
<< locali >>
rect 100 32 2536 128
<< locali >>
rect 93 25 157 135
<< m1 >>
rect 93 25 157 135
<< viali >>
rect 100 32 150 128
<< locali >>
rect 2479 25 2543 135
<< m1 >>
rect 2479 25 2543 135
<< viali >>
rect 2486 32 2536 128
<< labels >>
flabel m2 s 243 1982 386 2012 0 FreeSans 400 0 0 0 IN+
port 58 nsew signal bidirectional
flabel m2 s 819 2382 962 2412 0 FreeSans 400 0 0 0 IN-
port 59 nsew signal bidirectional
flabel locali s 0 8856 2636 8906 0 FreeSans 400 0 0 0 VDD
port 60 nsew signal bidirectional
flabel locali s 100 8756 2536 8806 0 FreeSans 400 0 0 0 VSS
port 61 nsew signal bidirectional
flabel m2 s 147 223 674 253 0 FreeSans 400 0 0 0 OUT
port 62 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1745590424
<< checkpaint >>
rect 0 0 1 1
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 1300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP diff1_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 1700
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 1300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP diff1_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 1700
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 3300
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 3700
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 3300
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 3700
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2500
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2260
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2500
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2260
box 0 0 832 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror2_MN4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 260
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror2_MN3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 260
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 900
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 900
box 0 0 576 400
use JNWATR_PCH_12C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2900
box 0 0 832 400
use JNWATR_PCH_12C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2900
box 0 0 832 400
<< locali >>
rect 100 4050 2164 4100
<< locali >>
rect 100 100 2164 150
<< m1 >>
rect 100 150 150 4050
<< m1 >>
rect 2114 150 2164 4050
<< locali >>
rect 93 4043 157 4107
<< m1 >>
rect 93 4043 157 4107
<< viali >>
rect 100 4050 150 4100
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2107 4043 2171 4107
<< m1 >>
rect 2107 4043 2171 4107
<< viali >>
rect 2114 4050 2164 4100
<< locali >>
rect 2107 93 2171 157
<< m1 >>
rect 2107 93 2171 157
<< viali >>
rect 2114 100 2164 150
<< locali >>
rect 0 4150 2264 4200
<< locali >>
rect 0 0 2264 50
<< m1 >>
rect 0 50 50 4150
<< m1 >>
rect 2214 50 2264 4150
<< locali >>
rect -7 4143 57 4207
<< m1 >>
rect -7 4143 57 4207
<< viali >>
rect 0 4150 50 4200
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2207 4143 2271 4207
<< m1 >>
rect 2207 4143 2271 4207
<< viali >>
rect 2214 4150 2264 4200
<< locali >>
rect 2207 -7 2271 57
<< m1 >>
rect 2207 -7 2271 57
<< viali >>
rect 2214 0 2264 50
<< locali >>
rect 1084 3600 1372 3640
<< locali >>
rect 1724 3480 1884 3520
<< locali >>
rect 252 3600 540 3640
<< locali >>
rect 1084 2800 1372 2840
<< locali >>
rect 252 2800 540 2840
<< locali >>
rect 892 2680 1052 2720
<< locali >>
rect 508 800 796 840
<< locali >>
rect 1084 800 1372 840
<< locali >>
rect 1468 680 1628 720
<< locali >>
rect 1084 1200 1372 1240
<< locali >>
rect 1468 1080 1628 1120
<< locali >>
rect 508 1200 796 1240
<< locali >>
rect 252 3200 540 3240
<< locali >>
rect 1084 3200 1372 3240
<< locali >>
rect 0 1772 2264 1868
<< locali >>
rect -7 1765 57 1875
<< m1 >>
rect -7 1765 57 1875
<< viali >>
rect 0 1772 50 1868
<< locali >>
rect 2207 1765 2271 1875
<< m1 >>
rect 2207 1765 2271 1875
<< viali >>
rect 2214 1772 2264 1868
<< locali >>
rect 100 3772 2164 3868
<< locali >>
rect 93 3765 157 3875
<< m1 >>
rect 93 3765 157 3875
<< viali >>
rect 100 3772 150 3868
<< locali >>
rect 2107 3765 2171 3875
<< m1 >>
rect 2107 3765 2171 3875
<< viali >>
rect 2114 3772 2164 3868
<< locali >>
rect 100 2332 2164 2428
<< locali >>
rect 93 2325 157 2435
<< m1 >>
rect 93 2325 157 2435
<< viali >>
rect 100 2332 150 2428
<< locali >>
rect 2107 2325 2171 2435
<< m1 >>
rect 2107 2325 2171 2435
<< viali >>
rect 2114 2332 2164 2428
<< locali >>
rect 0 332 2264 428
<< locali >>
rect -7 325 57 435
<< m1 >>
rect -7 325 57 435
<< viali >>
rect 0 332 50 428
<< locali >>
rect 2207 325 2271 435
<< m1 >>
rect 2207 325 2271 435
<< viali >>
rect 2214 332 2264 428
use COMP2 U1_COMP2 
transform 1 0 2314 0 1 0
box 0 0 1802 4250
use COMP2 U2_COMP2 
transform 1 0 0 0 1 5000
box 0 0 1802 4250
use COMP3 U3_COMP3 
transform 1 0 3604 0 1 5000
box 0 0 1802 4250
<< labels >>
flabel locali s 0 4150 2264 4200 0 FreeSans 400 0 0 0 VSS
port 118 nsew signal bidirectional
flabel locali s 100 4050 2164 4100 0 FreeSans 400 0 0 0 VDD
port 119 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1744043309
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 2000
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 1760
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 2000
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 1760
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 0
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 -240
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 -240
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 800
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 1200
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 800
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 1200
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 2800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 3200
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 2800
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 3200
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 2400
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 2400
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 576 0 1 400
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 0 0 1 400
box 0 0 576 400
<< locali >>
rect -250 3550 1402 3650
<< locali >>
rect -250 -450 1402 -350
<< m1 >>
rect -250 -350 -150 3550
<< m1 >>
rect 1302 -350 1402 3550
<< locali >>
rect -257 3543 -143 3657
<< m1 >>
rect -257 3543 -143 3657
<< viali >>
rect -250 3550 -150 3650
<< locali >>
rect -257 -457 -143 -343
<< m1 >>
rect -257 -457 -143 -343
<< viali >>
rect -250 -450 -150 -350
<< locali >>
rect 1295 3543 1409 3657
<< m1 >>
rect 1295 3543 1409 3657
<< viali >>
rect 1302 3550 1402 3650
<< locali >>
rect 1295 -457 1409 -343
<< m1 >>
rect 1295 -457 1409 -343
<< viali >>
rect 1302 -450 1402 -350
<< locali >>
rect -400 3700 1552 3800
<< locali >>
rect -400 -600 1552 -500
<< m1 >>
rect -400 -500 -300 3700
<< m1 >>
rect 1452 -500 1552 3700
<< locali >>
rect -407 3693 -293 3807
<< m1 >>
rect -407 3693 -293 3807
<< viali >>
rect -400 3700 -300 3800
<< locali >>
rect -407 -607 -293 -493
<< m1 >>
rect -407 -607 -293 -493
<< viali >>
rect -400 -600 -300 -500
<< locali >>
rect 1445 3693 1559 3807
<< m1 >>
rect 1445 3693 1559 3807
<< viali >>
rect 1452 3700 1552 3800
<< locali >>
rect 1445 -607 1559 -493
<< m1 >>
rect 1445 -607 1559 -493
<< viali >>
rect 1452 -600 1552 -500
<< locali >>
rect 528 300 816 340
<< locali >>
rect 912 180 1072 220
<< locali >>
rect -48 300 240 340
<< locali >>
rect -48 1100 240 1140
<< locali >>
rect 528 1100 816 1140
<< locali >>
rect 912 980 1072 1020
<< locali >>
rect -48 3100 240 3140
<< locali >>
rect 528 3100 816 3140
<< locali >>
rect 912 2980 1072 3020
<< locali >>
rect 528 2700 816 2740
<< locali >>
rect 912 2580 1072 2620
<< locali >>
rect -48 2700 240 2740
<< locali >>
rect 528 700 816 740
<< locali >>
rect -48 700 240 740
<< locali >>
rect -400 1832 1552 1928
<< locali >>
rect -407 1825 -293 1935
<< m1 >>
rect -407 1825 -293 1935
<< viali >>
rect -400 1832 -300 1928
<< locali >>
rect 1445 1825 1559 1935
<< m1 >>
rect 1445 1825 1559 1935
<< viali >>
rect 1452 1832 1552 1928
<< locali >>
rect -250 -168 1402 -72
<< locali >>
rect -257 -175 -143 -65
<< m1 >>
rect -257 -175 -143 -65
<< viali >>
rect -250 -168 -150 -72
<< locali >>
rect 1295 -175 1409 -65
<< m1 >>
rect 1295 -175 1409 -65
<< viali >>
rect 1302 -168 1402 -72
<< locali >>
rect -250 1272 1402 1368
<< locali >>
rect -257 1265 -143 1375
<< m1 >>
rect -257 1265 -143 1375
<< viali >>
rect -250 1272 -150 1368
<< locali >>
rect 1295 1265 1409 1375
<< m1 >>
rect 1295 1265 1409 1375
<< viali >>
rect 1302 1272 1402 1368
<< locali >>
rect -400 3272 1552 3368
<< locali >>
rect -407 3265 -293 3375
<< m1 >>
rect -407 3265 -293 3375
<< viali >>
rect -400 3272 -300 3368
<< locali >>
rect 1445 3265 1559 3375
<< m1 >>
rect 1445 3265 1559 3375
<< viali >>
rect 1452 3272 1552 3368
<< labels >>
flabel locali s -400 3700 1552 3800 0 FreeSans 400 0 0 0 VSS
port 47 nsew signal bidirectional
flabel locali s -250 3550 1402 3650 0 FreeSans 400 0 0 0 VDD
port 48 nsew signal bidirectional
<< properties >>
<< end >>
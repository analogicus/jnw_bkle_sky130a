magic
tech sky130A
magscale 1 1
timestamp 1745057841
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2260
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 2260
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 1300
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 1700
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 1300
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 1700
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 500
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 260
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 500
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 260
box 0 0 832 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 3300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 3700
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 3300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror2_MN3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 3700
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 2900
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 556 0 1 2900
box 0 0 576 400
use JNWATR_PCH_12C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1132 0 1 900
box 0 0 832 400
use JNWATR_PCH_12C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 900
box 0 0 832 400
<< locali >>
rect 100 4050 2164 4100
<< locali >>
rect 100 100 2164 150
<< m1 >>
rect 100 150 150 4050
<< m1 >>
rect 2114 150 2164 4050
<< locali >>
rect 93 4043 157 4107
<< m1 >>
rect 93 4043 157 4107
<< viali >>
rect 100 4050 150 4100
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2107 4043 2171 4107
<< m1 >>
rect 2107 4043 2171 4107
<< viali >>
rect 2114 4050 2164 4100
<< locali >>
rect 2107 93 2171 157
<< m1 >>
rect 2107 93 2171 157
<< viali >>
rect 2114 100 2164 150
<< locali >>
rect 0 4150 2264 4200
<< locali >>
rect 0 0 2264 50
<< m1 >>
rect 0 50 50 4150
<< m1 >>
rect 2214 50 2264 4150
<< locali >>
rect -7 4143 57 4207
<< m1 >>
rect -7 4143 57 4207
<< viali >>
rect 0 4150 50 4200
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2207 4143 2271 4207
<< m1 >>
rect 2207 4143 2271 4207
<< viali >>
rect 2214 4150 2264 4200
<< locali >>
rect 2207 -7 2271 57
<< m1 >>
rect 2207 -7 2271 57
<< viali >>
rect 2214 0 2264 50
<< locali >>
rect 1084 1600 1372 1640
<< locali >>
rect 1724 1480 1884 1520
<< locali >>
rect 252 1600 540 1640
<< locali >>
rect 252 800 540 840
<< locali >>
rect 1084 800 1372 840
<< locali >>
rect 1724 680 1884 720
<< locali >>
rect 508 3600 796 3640
<< locali >>
rect 1084 3600 1372 3640
<< locali >>
rect 1468 3480 1628 3520
<< locali >>
rect 1084 3200 1372 3240
<< locali >>
rect 1468 3080 1628 3120
<< locali >>
rect 508 3200 796 3240
<< locali >>
rect 1084 1200 1372 1240
<< locali >>
rect 252 1200 540 1240
<< locali >>
rect 0 2332 2264 2428
<< locali >>
rect -7 2325 57 2435
<< m1 >>
rect -7 2325 57 2435
<< viali >>
rect 0 2332 50 2428
<< locali >>
rect 2207 2325 2271 2435
<< m1 >>
rect 2207 2325 2271 2435
<< viali >>
rect 2214 2332 2264 2428
<< locali >>
rect 100 1772 2164 1868
<< locali >>
rect 93 1765 157 1875
<< m1 >>
rect 93 1765 157 1875
<< viali >>
rect 100 1772 150 1868
<< locali >>
rect 2107 1765 2171 1875
<< m1 >>
rect 2107 1765 2171 1875
<< viali >>
rect 2114 1772 2164 1868
<< locali >>
rect 100 332 2164 428
<< locali >>
rect 93 325 157 435
<< m1 >>
rect 93 325 157 435
<< viali >>
rect 100 332 150 428
<< locali >>
rect 2107 325 2171 435
<< m1 >>
rect 2107 325 2171 435
<< viali >>
rect 2114 332 2164 428
<< locali >>
rect 0 3772 2264 3868
<< locali >>
rect -7 3765 57 3875
<< m1 >>
rect -7 3765 57 3875
<< viali >>
rect 0 3772 50 3868
<< locali >>
rect 2207 3765 2271 3875
<< m1 >>
rect 2207 3765 2271 3875
<< viali >>
rect 2214 3772 2264 3868
use COMP2 U3_COMP2 
transform 1 0 2314 0 1 0
box 0 0 1802 4250
<< labels >>
flabel locali s 0 4150 2264 4200 0 FreeSans 400 0 0 0 VSS
port 6 nsew signal bidirectional
flabel locali s 100 4050 2164 4100 0 FreeSans 400 0 0 0 VDD
port 7 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1728915661
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 x1 ../JNW_ATR_SKY130A
transform 1 0 2500 0 1 1500
box 0 0 832 400
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform 1 0 4000 0 1 1500
box 0 0 512 400
use JNWTR_CAPX1 x4 ../JNW_TR_SKY130A
transform 1 0 5500 0 1 1500
box 0 0 540 540
use JNWTR_RES2 x3 ../JNW_TR_SKY130A
transform 1 0 7000 0 1 1500
box 0 0 324 1320
use JNWATR_NCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 1 0 8500 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x3 ../JNW_ATR_SKY130A
transform 1 0 10000 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x7 ../JNW_ATR_SKY130A
transform 1 0 11500 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x9 ../JNW_ATR_SKY130A
transform 1 0 13000 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x8 ../JNW_ATR_SKY130A
transform 1 0 14500 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x5 ../JNW_ATR_SKY130A
transform 1 0 16000 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform 1 0 17500 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 19000 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x10 ../JNW_ATR_SKY130A
transform 1 0 20500 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 x11 ../JNW_ATR_SKY130A
transform 1 0 22000 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x12 ../JNW_ATR_SKY130A
transform 1 0 23500 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 x13 ../JNW_ATR_SKY130A
transform 1 0 25000 0 1 1500
box 0 0 576 400
<< labels >>
<< properties >>
<< end >>
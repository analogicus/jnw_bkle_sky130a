magic
tech sky130A
magscale 1 1
timestamp 1729504246
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 x1 ../JNW_ATR_SKY130A
transform -1 0 99512 0 -1 940
box 0 0 832 400
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform -1 0 99192 0 -1 540
box 0 0 512 400
use JNWTR_CAPX1 x4 ../JNW_TR_SKY130A
transform -1 0 98680 0 -1 540
box 0 0 540 540
use JNWTR_RES2 x3 ../JNW_TR_SKY130A
transform 0 1 100000 -1 0 1264
box 0 0 324 1320
use JNWATR_NCH_4C5F0 x5 ../JNW_ATR_SKY130A
transform 0 -1 98280 1 0 2492
box 0 0 576 400
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform -1 0 98680 0 -1 1340
box 0 0 576 400
use JNWATR_PCH_4C5F0 x7 ../JNW_ATR_SKY130A
transform 1 0 98680 0 1 98680
box 0 0 576 400
use JNWATR_PCH_4C5F0 x8 ../JNW_ATR_SKY130A
transform 0 -1 98680 1 0 2492
box 0 0 576 400
use JNWATR_PCH_4C5F0 x9 ../JNW_ATR_SKY130A
transform 0 1 98280 -1 0 1916
box 0 0 576 400
use JNWATR_PCH_4C5F0 x10 ../JNW_ATR_SKY130A
transform 0 1 97880 -1 0 2492
box 0 0 576 400
use JNWATR_NCH_4C5F0 x11 ../JNW_ATR_SKY130A
transform 1 0 97480 0 1 97480
box 0 0 576 400
use JNWATR_NCH_4C5F0 x12 ../JNW_ATR_SKY130A
transform 0 1 97480 -1 0 1916
box 0 0 576 400
use JNWATR_NCH_4C5F0 x13 ../JNW_ATR_SKY130A
transform -1 0 97480 0 -1 1340
box 0 0 576 400
use JNWATR_NCH_4C5F0 x14 ../JNW_ATR_SKY130A
transform 0 -1 97880 1 0 1916
box 0 0 576 400
use JNWATR_PCH_4C5F0 x15 ../JNW_ATR_SKY130A
transform 1 0 98680 0 1 98680
box 0 0 576 400
use JNWATR_PCH_4C5F0 x16 ../JNW_ATR_SKY130A
transform 0 1 98680 -1 0 1916
box 0 0 576 400
<< labels >>
<< properties >>
<< end >>

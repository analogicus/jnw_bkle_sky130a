magic
tech sky130A
magscale 1 1
timestamp 1745918167
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5120
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWTR_CAPX1 None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4420
box 0 0 540 540
use JNWATR_PCH_4C5F0 None_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<9> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<8> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<7> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<6> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<5> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<4> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN1<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5360
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 5760
box 0 0 576 240
use JNWTR_RPPO8 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2300
box 0 0 1372 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 940 1720
use AALMISC_PNP_W3p40L3p40 load1_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6160
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<0> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 970 0 1 6160
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<1> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 970 0 1 7500
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<2> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 7500
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<3> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 970 0 1 8170
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<4> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 8170
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<5> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 970 0 1 6830
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<6> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 300 0 1 6830
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<7> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 970 0 1 8840
box 0 0 670 670
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< m3 >>
rect 373 5533 419 5587
<< via2 >>
rect 380 5540 412 5580
<< via1 >>
rect 380 5540 412 5580
<< m3 >>
rect 375 5237 405 5556
<< m2 >>
rect 375 5237 581 5267
<< m3 >>
rect 551 4436 581 5267
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m1 >>
rect 373 5533 419 5587
<< m2 >>
rect 373 5533 419 5587
<< via1 >>
rect 380 5540 412 5580
<< m2 >>
rect 368 5230 412 5274
<< m3 >>
rect 368 5230 412 5274
<< via2 >>
rect 375 5237 405 5267
<< m2 >>
rect 544 5230 588 5274
<< m3 >>
rect 544 5230 588 5274
<< via2 >>
rect 551 5237 581 5267
<< locali >>
rect 100 9860 1872 9910
<< locali >>
rect 100 100 1872 150
<< m1 >>
rect 100 150 150 9860
<< m1 >>
rect 1822 150 1872 9860
<< locali >>
rect 93 9853 157 9917
<< m1 >>
rect 93 9853 157 9917
<< viali >>
rect 100 9860 150 9910
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1815 9853 1879 9917
<< m1 >>
rect 1815 9853 1879 9917
<< viali >>
rect 1822 9860 1872 9910
<< locali >>
rect 1815 93 1879 157
<< m1 >>
rect 1815 93 1879 157
<< viali >>
rect 1822 100 1872 150
<< locali >>
rect 0 9960 1972 10010
<< locali >>
rect 0 0 1972 50
<< m1 >>
rect 0 50 50 9960
<< m1 >>
rect 1922 50 1972 9960
<< locali >>
rect -7 9953 57 10017
<< m1 >>
rect -7 9953 57 10017
<< viali >>
rect 0 9960 50 10010
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1915 9953 1979 10017
<< m1 >>
rect 1915 9953 1979 10017
<< viali >>
rect 1922 9960 1972 10010
<< locali >>
rect 1915 -7 1979 57
<< m1 >>
rect 1915 -7 1979 57
<< viali >>
rect 1922 0 1972 50
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 636 5540 796 5580
<< locali >>
rect 252 5660 540 5700
<< locali >>
rect 100 5192 1872 5288
<< locali >>
rect 93 5185 157 5295
<< m1 >>
rect 93 5185 157 5295
<< viali >>
rect 100 5192 150 5288
<< locali >>
rect 1815 5185 1879 5295
<< m1 >>
rect 1815 5185 1879 5295
<< viali >>
rect 1822 5192 1872 5288
<< locali >>
rect 0 3964 1972 4020
<< locali >>
rect -7 3957 57 4027
<< m1 >>
rect -7 3957 57 4027
<< viali >>
rect 0 3964 50 4020
<< locali >>
rect 1915 3957 1979 4027
<< m1 >>
rect 1915 3957 1979 4027
<< viali >>
rect 1922 3964 1972 4020
<< locali >>
rect 0 2300 1972 2356
<< locali >>
rect -7 2293 57 2363
<< m1 >>
rect -7 2293 57 2363
<< viali >>
rect 0 2300 50 2356
<< locali >>
rect 1915 2293 1979 2363
<< m1 >>
rect 1915 2293 1979 2363
<< viali >>
rect 1922 2300 1972 2356
<< locali >>
rect 0 2164 1972 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 1915 2157 1979 2227
<< m1 >>
rect 1915 2157 1979 2227
<< viali >>
rect 1922 2164 1972 2220
<< locali >>
rect 0 500 1972 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 1915 493 1979 563
<< m1 >>
rect 1915 493 1979 563
<< viali >>
rect 1922 500 1972 556
use OTA U1_OTA 
transform 1 0 2022 0 1 0
box 0 0 2886 10040
<< labels >>
flabel locali s 100 9860 1872 9910 0 FreeSans 400 0 0 0 VDD
port 35 nsew signal bidirectional
flabel locali s 0 9960 1972 10010 0 FreeSans 400 0 0 0 VSS
port 36 nsew signal bidirectional
flabel m1 s 636 5380 732 5420 0 FreeSans 400 0 0 0 OUT
port 37 nsew signal bidirectional
<< properties >>
<< end >>
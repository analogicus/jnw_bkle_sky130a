magic
tech sky130A
magscale 1 1
timestamp 1744381985
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_12C1F2 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 600
box 0 0 832 400
use JNWATR_NCH_12CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 1000
box 0 0 832 240
use JNWATR_NCH_12CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 400 0 1 360
box 0 0 832 240
<< locali >>
rect 150 1350 1482 1450
<< locali >>
rect 150 150 1482 250
<< m1 >>
rect 150 250 250 1350
<< m1 >>
rect 1382 250 1482 1350
<< locali >>
rect 143 1343 257 1457
<< m1 >>
rect 143 1343 257 1457
<< viali >>
rect 150 1350 250 1450
<< locali >>
rect 143 143 257 257
<< m1 >>
rect 143 143 257 257
<< viali >>
rect 150 150 250 250
<< locali >>
rect 1375 1343 1489 1457
<< m1 >>
rect 1375 1343 1489 1457
<< viali >>
rect 1382 1350 1482 1450
<< locali >>
rect 1375 143 1489 257
<< m1 >>
rect 1375 143 1489 257
<< viali >>
rect 1382 150 1482 250
<< locali >>
rect 0 1500 1632 1600
<< locali >>
rect 0 0 1632 100
<< m1 >>
rect 0 100 100 1500
<< m1 >>
rect 1532 100 1632 1500
<< locali >>
rect -7 1493 107 1607
<< m1 >>
rect -7 1493 107 1607
<< viali >>
rect 0 1500 100 1600
<< locali >>
rect -7 -7 107 107
<< m1 >>
rect -7 -7 107 107
<< viali >>
rect 0 0 100 100
<< locali >>
rect 1525 1493 1639 1607
<< m1 >>
rect 1525 1493 1639 1607
<< viali >>
rect 1532 1500 1632 1600
<< locali >>
rect 1525 -7 1639 107
<< m1 >>
rect 1525 -7 1639 107
<< viali >>
rect 1532 0 1632 100
<< locali >>
rect 352 900 640 940
<< locali >>
rect 992 780 1152 820
<< locali >>
rect 0 1072 1632 1168
<< locali >>
rect -7 1065 107 1175
<< m1 >>
rect -7 1065 107 1175
<< viali >>
rect 0 1072 100 1168
<< locali >>
rect 1525 1065 1639 1175
<< m1 >>
rect 1525 1065 1639 1175
<< viali >>
rect 1532 1072 1632 1168
<< locali >>
rect 0 432 1632 528
<< locali >>
rect -7 425 107 535
<< m1 >>
rect -7 425 107 535
<< viali >>
rect 0 432 100 528
<< locali >>
rect 1525 425 1639 535
<< m1 >>
rect 1525 425 1639 535
<< viali >>
rect 1532 432 1632 528
use COMP U1_COMP 
transform 1 0 1682 0 1 0
box 0 0 4306 2850
<< labels >>
flabel locali s 150 1350 1482 1450 0 FreeSans 400 0 0 0 VDD
port 4 nsew signal bidirectional
flabel locali s 0 1500 1632 1600 0 FreeSans 400 0 0 0 VSS
port 5 nsew signal bidirectional
<< properties >>
<< end >>
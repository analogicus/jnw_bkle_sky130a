magic
tech sky130A
magscale 1 1
timestamp 1745853979
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 7890
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP3<3>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8290
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 7890
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP3<2>_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 8290
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 7490
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 7490
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 7090
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 7090
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6690
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 6690
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6290
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 6050
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 6290
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 6050
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 9090
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 9490
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 8850
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9090
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9490
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8850
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2320
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 4170
box 0 0 2236 1720
<< m1 >>
rect 373 8063 419 8117
<< m2 >>
rect 373 8063 419 8117
<< m3 >>
rect 373 8063 419 8117
<< via2 >>
rect 380 8070 412 8110
<< via1 >>
rect 380 8070 412 8110
<< m1 >>
rect 949 8063 995 8117
<< m2 >>
rect 949 8063 995 8117
<< m3 >>
rect 949 8063 995 8117
<< via2 >>
rect 956 8070 988 8110
<< via1 >>
rect 956 8070 988 8110
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< m3 >>
rect 373 7663 419 7717
<< via2 >>
rect 380 7670 412 7710
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< m3 >>
rect 373 7663 419 7717
<< via2 >>
rect 380 7670 412 7710
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< m3 >>
rect 949 7663 995 7717
<< via2 >>
rect 956 7670 988 7710
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< m3 >>
rect 949 7663 995 7717
<< via2 >>
rect 956 7670 988 7710
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7263 995 7317
<< m2 >>
rect 949 7263 995 7317
<< m3 >>
rect 949 7263 995 7317
<< via2 >>
rect 956 7270 988 7310
<< via1 >>
rect 956 7270 988 7310
<< m1 >>
rect 373 6863 419 6917
<< m2 >>
rect 373 6863 419 6917
<< m3 >>
rect 373 6863 419 6917
<< via2 >>
rect 380 6870 412 6910
<< via1 >>
rect 380 6870 412 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< via1 >>
rect 956 6870 988 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< m3 >>
rect 949 6863 995 6917
<< via2 >>
rect 956 6870 988 6910
<< via1 >>
rect 956 6870 988 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< m3 >>
rect 949 6863 995 6917
<< via2 >>
rect 956 6870 988 6910
<< via1 >>
rect 956 6870 988 6910
<< m1 >>
rect 629 7103 739 7157
<< m2 >>
rect 629 7103 739 7157
<< m3 >>
rect 629 7103 739 7157
<< via2 >>
rect 636 7110 732 7150
<< via1 >>
rect 636 7110 732 7150
<< m1 >>
rect 1205 7103 1315 7157
<< m2 >>
rect 1205 7103 1315 7157
<< m3 >>
rect 1205 7103 1315 7157
<< via2 >>
rect 1212 7110 1308 7150
<< via1 >>
rect 1212 7110 1308 7150
<< m1 >>
rect 629 6703 739 6757
<< m2 >>
rect 629 6703 739 6757
<< m3 >>
rect 629 6703 739 6757
<< via2 >>
rect 636 6710 732 6750
<< via1 >>
rect 636 6710 732 6750
<< m1 >>
rect 629 6703 739 6757
<< m2 >>
rect 629 6703 739 6757
<< via1 >>
rect 636 6710 732 6750
<< m1 >>
rect 1205 6703 1315 6757
<< m2 >>
rect 1205 6703 1315 6757
<< via1 >>
rect 1212 6710 1308 6750
<< m1 >>
rect 1205 6703 1315 6757
<< m2 >>
rect 1205 6703 1315 6757
<< m3 >>
rect 1205 6703 1315 6757
<< via2 >>
rect 1212 6710 1308 6750
<< via1 >>
rect 1212 6710 1308 6750
<< m1 >>
rect 629 7903 739 7957
<< m2 >>
rect 629 7903 739 7957
<< m3 >>
rect 629 7903 739 7957
<< via2 >>
rect 636 7910 732 7950
<< via1 >>
rect 636 7910 732 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< m3 >>
rect 1205 7903 1315 7957
<< via2 >>
rect 1212 7910 1308 7950
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< m3 >>
rect 1205 7903 1315 7957
<< via2 >>
rect 1212 7910 1308 7950
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< m3 >>
rect 629 7503 739 7557
<< via2 >>
rect 636 7510 732 7550
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< m3 >>
rect 1205 7503 1315 7557
<< via2 >>
rect 1212 7510 1308 7550
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< m3 >>
rect 1205 7503 1315 7557
<< via2 >>
rect 1212 7510 1308 7550
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< m3 >>
rect 949 9263 995 9317
<< via2 >>
rect 956 9270 988 9310
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< m3 >>
rect 949 9263 995 9317
<< via2 >>
rect 956 9270 988 9310
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< m3 >>
rect 1205 9103 1315 9157
<< via2 >>
rect 1212 9110 1308 9150
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< m3 >>
rect 1205 9103 1315 9157
<< via2 >>
rect 1212 9110 1308 9150
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 373 9263 419 9317
<< m2 >>
rect 373 9263 419 9317
<< via1 >>
rect 380 9270 412 9310
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< m3 >>
rect 437 8183 547 8237
<< via2 >>
rect 444 8190 540 8230
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< m3 >>
rect 1013 8183 1123 8237
<< via2 >>
rect 1020 8190 1116 8230
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< m3 >>
rect 1013 8183 1123 8237
<< via2 >>
rect 1020 8190 1116 8230
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< m3 >>
rect 437 7783 547 7837
<< via2 >>
rect 444 7790 540 7830
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< m3 >>
rect 1013 7783 1123 7837
<< via2 >>
rect 1020 7790 1116 7830
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< m3 >>
rect 437 7383 547 7437
<< via2 >>
rect 444 7390 540 7430
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< m3 >>
rect 1013 7383 1123 7437
<< via2 >>
rect 1020 7390 1116 7430
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< m3 >>
rect 1013 7383 1123 7437
<< via2 >>
rect 1020 7390 1116 7430
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 437 6983 547 7037
<< m2 >>
rect 437 6983 547 7037
<< via1 >>
rect 444 6990 540 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< m3 >>
rect 1013 6983 1123 7037
<< via2 >>
rect 1020 6990 1116 7030
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< m3 >>
rect 629 6303 739 6357
<< via2 >>
rect 636 6310 732 6350
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 949 6463 995 6517
<< m2 >>
rect 949 6463 995 6517
<< m3 >>
rect 949 6463 995 6517
<< via2 >>
rect 956 6470 988 6510
<< via1 >>
rect 956 6470 988 6510
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< m3 >>
rect 1205 6303 1315 6357
<< via2 >>
rect 1212 6310 1308 6350
<< via1 >>
rect 1212 6310 1308 6350
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< m3 >>
rect 1205 6303 1315 6357
<< via2 >>
rect 1212 6310 1308 6350
<< via1 >>
rect 1212 6310 1308 6350
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< via1 >>
rect 1212 6310 1308 6350
<< locali >>
rect 2203 1953 2361 2087
<< m1 >>
rect 2203 1953 2361 2087
<< m2 >>
rect 2203 1953 2361 2087
<< via1 >>
rect 2210 1960 2354 2080
<< viali >>
rect 2210 1960 2354 2080
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< m2 >>
rect 475 1953 633 2087
<< m3 >>
rect 475 1953 633 2087
<< via2 >>
rect 482 1960 626 2080
<< via1 >>
rect 482 1960 626 2080
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< m2 >>
rect 2203 3773 2361 3907
<< via1 >>
rect 2210 3780 2354 3900
<< viali >>
rect 2210 3780 2354 3900
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< m2 >>
rect 475 3773 633 3907
<< m3 >>
rect 475 3773 633 3907
<< via2 >>
rect 482 3780 626 3900
<< via1 >>
rect 482 3780 626 3900
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< m2 >>
rect 2203 5623 2361 5757
<< via1 >>
rect 2210 5630 2354 5750
<< viali >>
rect 2210 5630 2354 5750
<< m3 >>
rect 954 7913 984 8088
<< m2 >>
rect 810 7913 984 7943
<< m3 >>
rect 810 7673 840 7943
<< m2 >>
rect 810 7673 984 7703
<< m3 >>
rect 954 7673 984 7703
<< m3 >>
rect 954 7513 984 7703
<< m2 >>
rect 810 7513 984 7543
<< m3 >>
rect 810 7289 840 7543
<< m2 >>
rect 522 7289 840 7319
<< m3 >>
rect 522 7145 552 7319
<< m2 >>
rect 234 7145 552 7175
<< m3 >>
rect 234 7145 264 7559
<< m2 >>
rect 234 7529 408 7559
<< m3 >>
rect 378 7529 408 7703
<< m3 >>
rect 378 7673 408 7703
<< m2 >>
rect 234 7673 408 7703
<< m3 >>
rect 234 7673 264 7959
<< m2 >>
rect 234 7929 408 7959
<< m3 >>
rect 378 7929 408 8088
<< m1 >>
rect 373 8063 419 8117
<< m2 >>
rect 373 8063 419 8117
<< via1 >>
rect 380 8070 412 8110
<< m1 >>
rect 949 8063 995 8117
<< m2 >>
rect 949 8063 995 8117
<< via1 >>
rect 956 8070 988 8110
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m2 >>
rect 947 7906 991 7950
<< m3 >>
rect 947 7906 991 7950
<< via2 >>
rect 954 7913 984 7943
<< m2 >>
rect 803 7906 847 7950
<< m3 >>
rect 803 7906 847 7950
<< via2 >>
rect 810 7913 840 7943
<< m2 >>
rect 803 7666 847 7710
<< m3 >>
rect 803 7666 847 7710
<< via2 >>
rect 810 7673 840 7703
<< m2 >>
rect 947 7666 991 7710
<< m3 >>
rect 947 7666 991 7710
<< via2 >>
rect 954 7673 984 7703
<< m2 >>
rect 947 7506 991 7550
<< m3 >>
rect 947 7506 991 7550
<< via2 >>
rect 954 7513 984 7543
<< m2 >>
rect 803 7506 847 7550
<< m3 >>
rect 803 7506 847 7550
<< via2 >>
rect 810 7513 840 7543
<< m2 >>
rect 803 7282 847 7326
<< m3 >>
rect 803 7282 847 7326
<< via2 >>
rect 810 7289 840 7319
<< m2 >>
rect 515 7282 559 7326
<< m3 >>
rect 515 7282 559 7326
<< via2 >>
rect 522 7289 552 7319
<< m2 >>
rect 515 7138 559 7182
<< m3 >>
rect 515 7138 559 7182
<< via2 >>
rect 522 7145 552 7175
<< m2 >>
rect 227 7138 271 7182
<< m3 >>
rect 227 7138 271 7182
<< via2 >>
rect 234 7145 264 7175
<< m2 >>
rect 227 7522 271 7566
<< m3 >>
rect 227 7522 271 7566
<< via2 >>
rect 234 7529 264 7559
<< m2 >>
rect 371 7522 415 7566
<< m3 >>
rect 371 7522 415 7566
<< via2 >>
rect 378 7529 408 7559
<< m2 >>
rect 371 7666 415 7710
<< m3 >>
rect 371 7666 415 7710
<< via2 >>
rect 378 7673 408 7703
<< m2 >>
rect 227 7666 271 7710
<< m3 >>
rect 227 7666 271 7710
<< via2 >>
rect 234 7673 264 7703
<< m2 >>
rect 227 7922 271 7966
<< m3 >>
rect 227 7922 271 7966
<< via2 >>
rect 234 7929 264 7959
<< m2 >>
rect 371 7922 415 7966
<< m3 >>
rect 371 7922 415 7966
<< via2 >>
rect 378 7929 408 7959
<< m3 >>
rect 954 7113 984 7288
<< m2 >>
rect 810 7113 984 7143
<< m3 >>
rect 810 6873 840 7143
<< m2 >>
rect 810 6873 984 6903
<< m3 >>
rect 954 6873 984 6903
<< m3 >>
rect 954 6681 984 6903
<< m2 >>
rect 810 6681 984 6711
<< m3 >>
rect 810 6521 840 6711
<< m2 >>
rect 522 6521 840 6551
<< m3 >>
rect 522 6361 552 6551
<< m2 >>
rect 234 6361 552 6391
<< m3 >>
rect 234 6361 264 6743
<< m2 >>
rect 234 6713 408 6743
<< m3 >>
rect 378 6713 408 6888
<< m1 >>
rect 949 7263 995 7317
<< m2 >>
rect 949 7263 995 7317
<< via1 >>
rect 956 7270 988 7310
<< m1 >>
rect 373 6863 419 6917
<< m2 >>
rect 373 6863 419 6917
<< via1 >>
rect 380 6870 412 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< via1 >>
rect 956 6870 988 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< via1 >>
rect 956 6870 988 6910
<< m1 >>
rect 949 6863 995 6917
<< m2 >>
rect 949 6863 995 6917
<< via1 >>
rect 956 6870 988 6910
<< m2 >>
rect 947 7106 991 7150
<< m3 >>
rect 947 7106 991 7150
<< via2 >>
rect 954 7113 984 7143
<< m2 >>
rect 803 7106 847 7150
<< m3 >>
rect 803 7106 847 7150
<< via2 >>
rect 810 7113 840 7143
<< m2 >>
rect 803 6866 847 6910
<< m3 >>
rect 803 6866 847 6910
<< via2 >>
rect 810 6873 840 6903
<< m2 >>
rect 947 6866 991 6910
<< m3 >>
rect 947 6866 991 6910
<< via2 >>
rect 954 6873 984 6903
<< m2 >>
rect 947 6674 991 6718
<< m3 >>
rect 947 6674 991 6718
<< via2 >>
rect 954 6681 984 6711
<< m2 >>
rect 803 6674 847 6718
<< m3 >>
rect 803 6674 847 6718
<< via2 >>
rect 810 6681 840 6711
<< m2 >>
rect 803 6514 847 6558
<< m3 >>
rect 803 6514 847 6558
<< via2 >>
rect 810 6521 840 6551
<< m2 >>
rect 515 6514 559 6558
<< m3 >>
rect 515 6514 559 6558
<< via2 >>
rect 522 6521 552 6551
<< m2 >>
rect 515 6354 559 6398
<< m3 >>
rect 515 6354 559 6398
<< via2 >>
rect 522 6361 552 6391
<< m2 >>
rect 227 6354 271 6398
<< m3 >>
rect 227 6354 271 6398
<< via2 >>
rect 234 6361 264 6391
<< m2 >>
rect 227 6706 271 6750
<< m3 >>
rect 227 6706 271 6750
<< via2 >>
rect 234 6713 264 6743
<< m2 >>
rect 371 6706 415 6750
<< m3 >>
rect 371 6706 415 6750
<< via2 >>
rect 378 6713 408 6743
<< m3 >>
rect 667 6713 697 7128
<< m2 >>
rect 667 6713 1273 6743
<< m3 >>
rect 1243 6713 1273 7128
<< m1 >>
rect 629 7103 739 7157
<< m2 >>
rect 629 7103 739 7157
<< via1 >>
rect 636 7110 732 7150
<< m1 >>
rect 1205 7103 1315 7157
<< m2 >>
rect 1205 7103 1315 7157
<< via1 >>
rect 1212 7110 1308 7150
<< m1 >>
rect 629 6703 739 6757
<< m2 >>
rect 629 6703 739 6757
<< via1 >>
rect 636 6710 732 6750
<< m1 >>
rect 629 6703 739 6757
<< m2 >>
rect 629 6703 739 6757
<< via1 >>
rect 636 6710 732 6750
<< m1 >>
rect 1205 6703 1315 6757
<< m2 >>
rect 1205 6703 1315 6757
<< via1 >>
rect 1212 6710 1308 6750
<< m1 >>
rect 1205 6703 1315 6757
<< m2 >>
rect 1205 6703 1315 6757
<< via1 >>
rect 1212 6710 1308 6750
<< m2 >>
rect 660 6706 704 6750
<< m3 >>
rect 660 6706 704 6750
<< via2 >>
rect 667 6713 697 6743
<< m2 >>
rect 1236 6706 1280 6750
<< m3 >>
rect 1236 6706 1280 6750
<< via2 >>
rect 1243 6713 1273 6743
<< m2 >>
rect 394 9274 985 9304
<< m3 >>
rect 955 9274 985 9304
<< m3 >>
rect 955 9114 985 9304
<< m2 >>
rect 955 9114 1273 9144
<< m3 >>
rect 1243 9114 1273 9144
<< m3 >>
rect 1243 7914 1273 9144
<< m3 >>
rect 1243 7914 1273 7944
<< m2 >>
rect 1243 7914 1417 7944
<< m3 >>
rect 1387 7658 1417 7944
<< m2 >>
rect 1243 7658 1417 7688
<< m3 >>
rect 1243 7514 1273 7688
<< m3 >>
rect 1243 7514 1273 7544
<< m2 >>
rect 1243 7514 1513 7544
<< m3 >>
rect 1483 7514 1513 8184
<< m2 >>
rect 1339 8154 1513 8184
<< m3 >>
rect 1339 8154 1369 8344
<< m2 >>
rect 811 8314 1369 8344
<< m3 >>
rect 811 8074 841 8344
<< m2 >>
rect 667 8074 841 8104
<< m3 >>
rect 667 7529 697 8104
<< m1 >>
rect 629 7903 739 7957
<< m2 >>
rect 629 7903 739 7957
<< via1 >>
rect 636 7910 732 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 373 9263 419 9317
<< m2 >>
rect 373 9263 419 9317
<< via1 >>
rect 380 9270 412 9310
<< m2 >>
rect 948 9267 992 9311
<< m3 >>
rect 948 9267 992 9311
<< via2 >>
rect 955 9274 985 9304
<< m2 >>
rect 948 9107 992 9151
<< m3 >>
rect 948 9107 992 9151
<< via2 >>
rect 955 9114 985 9144
<< m2 >>
rect 1236 9107 1280 9151
<< m3 >>
rect 1236 9107 1280 9151
<< via2 >>
rect 1243 9114 1273 9144
<< m2 >>
rect 1236 7907 1280 7951
<< m3 >>
rect 1236 7907 1280 7951
<< via2 >>
rect 1243 7914 1273 7944
<< m2 >>
rect 1380 7907 1424 7951
<< m3 >>
rect 1380 7907 1424 7951
<< via2 >>
rect 1387 7914 1417 7944
<< m2 >>
rect 1380 7651 1424 7695
<< m3 >>
rect 1380 7651 1424 7695
<< via2 >>
rect 1387 7658 1417 7688
<< m2 >>
rect 1236 7651 1280 7695
<< m3 >>
rect 1236 7651 1280 7695
<< via2 >>
rect 1243 7658 1273 7688
<< m2 >>
rect 1236 7507 1280 7551
<< m3 >>
rect 1236 7507 1280 7551
<< via2 >>
rect 1243 7514 1273 7544
<< m2 >>
rect 1476 7507 1520 7551
<< m3 >>
rect 1476 7507 1520 7551
<< via2 >>
rect 1483 7514 1513 7544
<< m2 >>
rect 1476 8147 1520 8191
<< m3 >>
rect 1476 8147 1520 8191
<< via2 >>
rect 1483 8154 1513 8184
<< m2 >>
rect 1332 8147 1376 8191
<< m3 >>
rect 1332 8147 1376 8191
<< via2 >>
rect 1339 8154 1369 8184
<< m2 >>
rect 1332 8307 1376 8351
<< m3 >>
rect 1332 8307 1376 8351
<< via2 >>
rect 1339 8314 1369 8344
<< m2 >>
rect 804 8307 848 8351
<< m3 >>
rect 804 8307 848 8351
<< via2 >>
rect 811 8314 841 8344
<< m2 >>
rect 804 8067 848 8111
<< m3 >>
rect 804 8067 848 8111
<< via2 >>
rect 811 8074 841 8104
<< m2 >>
rect 660 8067 704 8111
<< m3 >>
rect 660 8067 704 8111
<< via2 >>
rect 667 8074 697 8104
<< m3 >>
rect 668 6163 698 6322
<< m2 >>
rect 140 6163 698 6193
<< m3 >>
rect 140 6163 170 7025
<< m2 >>
rect 140 6995 506 7025
<< m2 >>
rect 668 6307 1098 6337
<< m3 >>
rect 1068 6307 1098 6529
<< m2 >>
rect 1068 6499 1418 6529
<< m3 >>
rect 1388 6499 1418 7009
<< m2 >>
rect 1068 6979 1418 7009
<< m3 >>
rect 1068 6979 1098 7425
<< m2 >>
rect 476 7395 1098 7425
<< m3 >>
rect 476 7395 506 7425
<< m2 >>
rect 140 7395 506 7425
<< m3 >>
rect 140 7395 170 7825
<< m2 >>
rect 140 7795 506 7825
<< m3 >>
rect 476 7795 506 8225
<< m2 >>
rect 476 8195 1082 8225
<< m3 >>
rect 1052 8195 1082 8225
<< m3 >>
rect 1052 8195 1082 8433
<< m2 >>
rect 1052 8403 1610 8433
<< m3 >>
rect 1580 7795 1610 8433
<< m2 >>
rect 1052 7795 1610 7825
<< m3 >>
rect 1052 7395 1082 7825
<< m2 >>
rect 1052 7395 1418 7425
<< m3 >>
rect 1388 6995 1418 7425
<< m2 >>
rect 1067 6995 1418 7025
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 437 7383 547 7437
<< m2 >>
rect 437 7383 547 7437
<< via1 >>
rect 444 7390 540 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 1013 7383 1123 7437
<< m2 >>
rect 1013 7383 1123 7437
<< via1 >>
rect 1020 7390 1116 7430
<< m1 >>
rect 437 6983 547 7037
<< m2 >>
rect 437 6983 547 7037
<< via1 >>
rect 444 6990 540 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 1013 6983 1123 7037
<< m2 >>
rect 1013 6983 1123 7037
<< via1 >>
rect 1020 6990 1116 7030
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m2 >>
rect 661 6156 705 6200
<< m3 >>
rect 661 6156 705 6200
<< via2 >>
rect 668 6163 698 6193
<< m2 >>
rect 133 6156 177 6200
<< m3 >>
rect 133 6156 177 6200
<< via2 >>
rect 140 6163 170 6193
<< m2 >>
rect 133 6988 177 7032
<< m3 >>
rect 133 6988 177 7032
<< via2 >>
rect 140 6995 170 7025
<< m2 >>
rect 1061 6300 1105 6344
<< m3 >>
rect 1061 6300 1105 6344
<< via2 >>
rect 1068 6307 1098 6337
<< m2 >>
rect 1061 6492 1105 6536
<< m3 >>
rect 1061 6492 1105 6536
<< via2 >>
rect 1068 6499 1098 6529
<< m2 >>
rect 1381 6492 1425 6536
<< m3 >>
rect 1381 6492 1425 6536
<< via2 >>
rect 1388 6499 1418 6529
<< m2 >>
rect 1381 6972 1425 7016
<< m3 >>
rect 1381 6972 1425 7016
<< via2 >>
rect 1388 6979 1418 7009
<< m2 >>
rect 1061 6972 1105 7016
<< m3 >>
rect 1061 6972 1105 7016
<< via2 >>
rect 1068 6979 1098 7009
<< m2 >>
rect 1061 7388 1105 7432
<< m3 >>
rect 1061 7388 1105 7432
<< via2 >>
rect 1068 7395 1098 7425
<< m2 >>
rect 469 7388 513 7432
<< m3 >>
rect 469 7388 513 7432
<< via2 >>
rect 476 7395 506 7425
<< m2 >>
rect 469 7388 513 7432
<< m3 >>
rect 469 7388 513 7432
<< via2 >>
rect 476 7395 506 7425
<< m2 >>
rect 133 7388 177 7432
<< m3 >>
rect 133 7388 177 7432
<< via2 >>
rect 140 7395 170 7425
<< m2 >>
rect 133 7788 177 7832
<< m3 >>
rect 133 7788 177 7832
<< via2 >>
rect 140 7795 170 7825
<< m2 >>
rect 469 7788 513 7832
<< m3 >>
rect 469 7788 513 7832
<< via2 >>
rect 476 7795 506 7825
<< m2 >>
rect 469 8188 513 8232
<< m3 >>
rect 469 8188 513 8232
<< via2 >>
rect 476 8195 506 8225
<< m2 >>
rect 1045 8188 1089 8232
<< m3 >>
rect 1045 8188 1089 8232
<< via2 >>
rect 1052 8195 1082 8225
<< m2 >>
rect 1045 8396 1089 8440
<< m3 >>
rect 1045 8396 1089 8440
<< via2 >>
rect 1052 8403 1082 8433
<< m2 >>
rect 1573 8396 1617 8440
<< m3 >>
rect 1573 8396 1617 8440
<< via2 >>
rect 1580 8403 1610 8433
<< m2 >>
rect 1573 7788 1617 7832
<< m3 >>
rect 1573 7788 1617 7832
<< via2 >>
rect 1580 7795 1610 7825
<< m2 >>
rect 1045 7788 1089 7832
<< m3 >>
rect 1045 7788 1089 7832
<< via2 >>
rect 1052 7795 1082 7825
<< m2 >>
rect 1045 7388 1089 7432
<< m3 >>
rect 1045 7388 1089 7432
<< via2 >>
rect 1052 7395 1082 7425
<< m2 >>
rect 1381 7388 1425 7432
<< m3 >>
rect 1381 7388 1425 7432
<< via2 >>
rect 1388 7395 1418 7425
<< m2 >>
rect 1381 6988 1425 7032
<< m3 >>
rect 1381 6988 1425 7032
<< via2 >>
rect 1388 6995 1418 7025
<< m2 >>
rect 2105 2007 2280 2037
<< m3 >>
rect 2105 2007 2135 2293
<< m2 >>
rect 1929 2263 2135 2293
<< m3 >>
rect 1929 2263 1959 2757
<< m2 >>
rect 1689 2727 1959 2757
<< m3 >>
rect 1689 2727 1719 3925
<< m2 >>
rect 1529 3895 1719 3925
<< m3 >>
rect 1529 3895 1559 6005
<< m2 >>
rect 1385 5975 1559 6005
<< m3 >>
rect 1385 5975 1415 6149
<< m2 >>
rect 1241 6119 1415 6149
<< m3 >>
rect 1241 6119 1271 6341
<< m3 >>
rect 1241 6311 1271 6341
<< m2 >>
rect 1241 6311 1559 6341
<< m3 >>
rect 1529 6311 1559 6485
<< m2 >>
rect 1529 6455 1703 6485
<< m3 >>
rect 1673 6215 1703 6485
<< m2 >>
rect 953 6215 1703 6245
<< m3 >>
rect 953 6215 983 6486
<< m1 >>
rect 949 6463 995 6517
<< m2 >>
rect 949 6463 995 6517
<< via1 >>
rect 956 6470 988 6510
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< via1 >>
rect 1212 6310 1308 6350
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< via1 >>
rect 1212 6310 1308 6350
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< via1 >>
rect 1212 6310 1308 6350
<< locali >>
rect 2203 1953 2361 2087
<< m1 >>
rect 2203 1953 2361 2087
<< viali >>
rect 2210 1960 2354 2080
<< m2 >>
rect 2098 2000 2142 2044
<< m3 >>
rect 2098 2000 2142 2044
<< via2 >>
rect 2105 2007 2135 2037
<< m2 >>
rect 2098 2256 2142 2300
<< m3 >>
rect 2098 2256 2142 2300
<< via2 >>
rect 2105 2263 2135 2293
<< m2 >>
rect 1922 2256 1966 2300
<< m3 >>
rect 1922 2256 1966 2300
<< via2 >>
rect 1929 2263 1959 2293
<< m2 >>
rect 1922 2720 1966 2764
<< m3 >>
rect 1922 2720 1966 2764
<< via2 >>
rect 1929 2727 1959 2757
<< m2 >>
rect 1682 2720 1726 2764
<< m3 >>
rect 1682 2720 1726 2764
<< via2 >>
rect 1689 2727 1719 2757
<< m2 >>
rect 1682 3888 1726 3932
<< m3 >>
rect 1682 3888 1726 3932
<< via2 >>
rect 1689 3895 1719 3925
<< m2 >>
rect 1522 3888 1566 3932
<< m3 >>
rect 1522 3888 1566 3932
<< via2 >>
rect 1529 3895 1559 3925
<< m2 >>
rect 1522 5968 1566 6012
<< m3 >>
rect 1522 5968 1566 6012
<< via2 >>
rect 1529 5975 1559 6005
<< m2 >>
rect 1378 5968 1422 6012
<< m3 >>
rect 1378 5968 1422 6012
<< via2 >>
rect 1385 5975 1415 6005
<< m2 >>
rect 1378 6112 1422 6156
<< m3 >>
rect 1378 6112 1422 6156
<< via2 >>
rect 1385 6119 1415 6149
<< m2 >>
rect 1234 6112 1278 6156
<< m3 >>
rect 1234 6112 1278 6156
<< via2 >>
rect 1241 6119 1271 6149
<< m2 >>
rect 1234 6304 1278 6348
<< m3 >>
rect 1234 6304 1278 6348
<< via2 >>
rect 1241 6311 1271 6341
<< m2 >>
rect 1522 6304 1566 6348
<< m3 >>
rect 1522 6304 1566 6348
<< via2 >>
rect 1529 6311 1559 6341
<< m2 >>
rect 1522 6448 1566 6492
<< m3 >>
rect 1522 6448 1566 6492
<< via2 >>
rect 1529 6455 1559 6485
<< m2 >>
rect 1666 6448 1710 6492
<< m3 >>
rect 1666 6448 1710 6492
<< via2 >>
rect 1673 6455 1703 6485
<< m2 >>
rect 1666 6208 1710 6252
<< m3 >>
rect 1666 6208 1710 6252
<< via2 >>
rect 1673 6215 1703 6245
<< m2 >>
rect 946 6208 990 6252
<< m3 >>
rect 946 6208 990 6252
<< via2 >>
rect 953 6215 983 6245
<< m3 >>
rect 534 2018 564 2193
<< m2 >>
rect 534 2163 772 2193
<< m3 >>
rect 742 2163 772 2385
<< m2 >>
rect 742 2355 916 2385
<< m3 >>
rect 886 2355 916 2545
<< m2 >>
rect 886 2515 1060 2545
<< m3 >>
rect 1030 2515 1060 2721
<< m2 >>
rect 1030 2691 1204 2721
<< m3 >>
rect 1174 2691 1204 2929
<< m2 >>
rect 1174 2899 1380 2929
<< m3 >>
rect 1350 2899 1380 3249
<< m2 >>
rect 1350 3219 1604 3249
<< m3 >>
rect 1574 3219 1604 3537
<< m2 >>
rect 1574 3507 1876 3537
<< m3 >>
rect 1846 3507 1876 3697
<< m2 >>
rect 1846 3667 2020 3697
<< m3 >>
rect 1990 3667 2020 3857
<< m2 >>
rect 1990 3827 2277 3857
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< viali >>
rect 2210 3780 2354 3900
<< m2 >>
rect 527 2156 571 2200
<< m3 >>
rect 527 2156 571 2200
<< via2 >>
rect 534 2163 564 2193
<< m2 >>
rect 735 2156 779 2200
<< m3 >>
rect 735 2156 779 2200
<< via2 >>
rect 742 2163 772 2193
<< m2 >>
rect 735 2348 779 2392
<< m3 >>
rect 735 2348 779 2392
<< via2 >>
rect 742 2355 772 2385
<< m2 >>
rect 879 2348 923 2392
<< m3 >>
rect 879 2348 923 2392
<< via2 >>
rect 886 2355 916 2385
<< m2 >>
rect 879 2508 923 2552
<< m3 >>
rect 879 2508 923 2552
<< via2 >>
rect 886 2515 916 2545
<< m2 >>
rect 1023 2508 1067 2552
<< m3 >>
rect 1023 2508 1067 2552
<< via2 >>
rect 1030 2515 1060 2545
<< m2 >>
rect 1023 2684 1067 2728
<< m3 >>
rect 1023 2684 1067 2728
<< via2 >>
rect 1030 2691 1060 2721
<< m2 >>
rect 1167 2684 1211 2728
<< m3 >>
rect 1167 2684 1211 2728
<< via2 >>
rect 1174 2691 1204 2721
<< m2 >>
rect 1167 2892 1211 2936
<< m3 >>
rect 1167 2892 1211 2936
<< via2 >>
rect 1174 2899 1204 2929
<< m2 >>
rect 1343 2892 1387 2936
<< m3 >>
rect 1343 2892 1387 2936
<< via2 >>
rect 1350 2899 1380 2929
<< m2 >>
rect 1343 3212 1387 3256
<< m3 >>
rect 1343 3212 1387 3256
<< via2 >>
rect 1350 3219 1380 3249
<< m2 >>
rect 1567 3212 1611 3256
<< m3 >>
rect 1567 3212 1611 3256
<< via2 >>
rect 1574 3219 1604 3249
<< m2 >>
rect 1567 3500 1611 3544
<< m3 >>
rect 1567 3500 1611 3544
<< via2 >>
rect 1574 3507 1604 3537
<< m2 >>
rect 1839 3500 1883 3544
<< m3 >>
rect 1839 3500 1883 3544
<< via2 >>
rect 1846 3507 1876 3537
<< m2 >>
rect 1839 3660 1883 3704
<< m3 >>
rect 1839 3660 1883 3704
<< via2 >>
rect 1846 3667 1876 3697
<< m2 >>
rect 1983 3660 2027 3704
<< m3 >>
rect 1983 3660 2027 3704
<< via2 >>
rect 1990 3667 2020 3697
<< m2 >>
rect 1983 3820 2027 3864
<< m3 >>
rect 1983 3820 2027 3864
<< via2 >>
rect 1990 3827 2020 3857
<< m3 >>
rect 534 3840 564 4095
<< m2 >>
rect 534 4065 740 4095
<< m3 >>
rect 710 4065 740 4271
<< m2 >>
rect 710 4241 980 4271
<< m3 >>
rect 950 4241 980 4447
<< m2 >>
rect 950 4417 1252 4447
<< m3 >>
rect 1222 4417 1252 4639
<< m2 >>
rect 1222 4609 1428 4639
<< m3 >>
rect 1398 4609 1428 4815
<< m2 >>
rect 1398 4785 1764 4815
<< m3 >>
rect 1734 4785 1764 5151
<< m2 >>
rect 1734 5121 1908 5151
<< m3 >>
rect 1878 5121 1908 5503
<< m2 >>
rect 1878 5473 2068 5503
<< m3 >>
rect 2038 5473 2068 5695
<< m2 >>
rect 2038 5665 2277 5695
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< viali >>
rect 2210 5630 2354 5750
<< m2 >>
rect 527 4058 571 4102
<< m3 >>
rect 527 4058 571 4102
<< via2 >>
rect 534 4065 564 4095
<< m2 >>
rect 703 4058 747 4102
<< m3 >>
rect 703 4058 747 4102
<< via2 >>
rect 710 4065 740 4095
<< m2 >>
rect 703 4234 747 4278
<< m3 >>
rect 703 4234 747 4278
<< via2 >>
rect 710 4241 740 4271
<< m2 >>
rect 943 4234 987 4278
<< m3 >>
rect 943 4234 987 4278
<< via2 >>
rect 950 4241 980 4271
<< m2 >>
rect 943 4410 987 4454
<< m3 >>
rect 943 4410 987 4454
<< via2 >>
rect 950 4417 980 4447
<< m2 >>
rect 1215 4410 1259 4454
<< m3 >>
rect 1215 4410 1259 4454
<< via2 >>
rect 1222 4417 1252 4447
<< m2 >>
rect 1215 4602 1259 4646
<< m3 >>
rect 1215 4602 1259 4646
<< via2 >>
rect 1222 4609 1252 4639
<< m2 >>
rect 1391 4602 1435 4646
<< m3 >>
rect 1391 4602 1435 4646
<< via2 >>
rect 1398 4609 1428 4639
<< m2 >>
rect 1391 4778 1435 4822
<< m3 >>
rect 1391 4778 1435 4822
<< via2 >>
rect 1398 4785 1428 4815
<< m2 >>
rect 1727 4778 1771 4822
<< m3 >>
rect 1727 4778 1771 4822
<< via2 >>
rect 1734 4785 1764 4815
<< m2 >>
rect 1727 5114 1771 5158
<< m3 >>
rect 1727 5114 1771 5158
<< via2 >>
rect 1734 5121 1764 5151
<< m2 >>
rect 1871 5114 1915 5158
<< m3 >>
rect 1871 5114 1915 5158
<< via2 >>
rect 1878 5121 1908 5151
<< m2 >>
rect 1871 5466 1915 5510
<< m3 >>
rect 1871 5466 1915 5510
<< via2 >>
rect 1878 5473 1908 5503
<< m2 >>
rect 2031 5466 2075 5510
<< m3 >>
rect 2031 5466 2075 5510
<< via2 >>
rect 2038 5473 2068 5503
<< m2 >>
rect 2031 5658 2075 5702
<< m3 >>
rect 2031 5658 2075 5702
<< via2 >>
rect 2038 5665 2068 5695
<< locali >>
rect 100 9840 2736 9890
<< locali >>
rect 100 100 2736 150
<< m1 >>
rect 100 150 150 9840
<< m1 >>
rect 2686 150 2736 9840
<< locali >>
rect 93 9833 157 9897
<< m1 >>
rect 93 9833 157 9897
<< viali >>
rect 100 9840 150 9890
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2679 9833 2743 9897
<< m1 >>
rect 2679 9833 2743 9897
<< viali >>
rect 2686 9840 2736 9890
<< locali >>
rect 2679 93 2743 157
<< m1 >>
rect 2679 93 2743 157
<< viali >>
rect 2686 100 2736 150
<< locali >>
rect 0 9940 2836 9990
<< locali >>
rect 0 0 2836 50
<< m1 >>
rect 0 50 50 9940
<< m1 >>
rect 2786 50 2836 9940
<< locali >>
rect -7 9933 57 9997
<< m1 >>
rect -7 9933 57 9997
<< viali >>
rect 0 9940 50 9990
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2779 9933 2843 9997
<< m1 >>
rect 2779 9933 2843 9997
<< viali >>
rect 2786 9940 2836 9990
<< locali >>
rect 2779 -7 2843 57
<< m1 >>
rect 2779 -7 2843 57
<< viali >>
rect 2786 0 2836 50
<< locali >>
rect 252 6590 540 6630
<< locali >>
rect 828 6590 1116 6630
<< locali >>
rect 1212 6470 1372 6510
<< locali >>
rect 828 9390 1116 9430
<< locali >>
rect 1212 9270 1372 9310
<< locali >>
rect 252 9390 540 9430
<< locali >>
rect 100 8362 2736 8458
<< locali >>
rect 93 8355 157 8465
<< m1 >>
rect 93 8355 157 8465
<< viali >>
rect 100 8362 150 8458
<< locali >>
rect 2679 8355 2743 8465
<< m1 >>
rect 2679 8355 2743 8465
<< viali >>
rect 2686 8362 2736 8458
<< locali >>
rect 100 6122 2736 6218
<< locali >>
rect 93 6115 157 6225
<< m1 >>
rect 93 6115 157 6225
<< viali >>
rect 100 6122 150 6218
<< locali >>
rect 2679 6115 2743 6225
<< m1 >>
rect 2679 6115 2743 6225
<< viali >>
rect 2686 6122 2736 6218
<< locali >>
rect 0 9562 2836 9658
<< locali >>
rect -7 9555 57 9665
<< m1 >>
rect -7 9555 57 9665
<< viali >>
rect 0 9562 50 9658
<< locali >>
rect 2779 9555 2843 9665
<< m1 >>
rect 2779 9555 2843 9665
<< viali >>
rect 2786 9562 2836 9658
<< locali >>
rect 0 8922 2836 9018
<< locali >>
rect -7 8915 57 9025
<< m1 >>
rect -7 8915 57 9025
<< viali >>
rect 0 8922 50 9018
<< locali >>
rect 2779 8915 2843 9025
<< m1 >>
rect 2779 8915 2843 9025
<< viali >>
rect 2786 8922 2836 9018
<< locali >>
rect 308 5630 626 5750
<< locali >>
rect 0 2164 2836 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 2779 2157 2843 2227
<< m1 >>
rect 2779 2157 2843 2227
<< viali >>
rect 2786 2164 2836 2220
<< locali >>
rect 0 500 2836 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 2779 493 2843 563
<< m1 >>
rect 2779 493 2843 563
<< viali >>
rect 2786 500 2836 556
<< locali >>
rect 0 3984 2836 4040
<< locali >>
rect -7 3977 57 4047
<< m1 >>
rect -7 3977 57 4047
<< viali >>
rect 0 3984 50 4040
<< locali >>
rect 2779 3977 2843 4047
<< m1 >>
rect 2779 3977 2843 4047
<< viali >>
rect 2786 3984 2836 4040
<< locali >>
rect 0 2320 2836 2376
<< locali >>
rect -7 2313 57 2383
<< m1 >>
rect -7 2313 57 2383
<< viali >>
rect 0 2320 50 2376
<< locali >>
rect 2779 2313 2843 2383
<< m1 >>
rect 2779 2313 2843 2383
<< viali >>
rect 2786 2320 2836 2376
<< locali >>
rect 0 5834 2836 5890
<< locali >>
rect -7 5827 57 5897
<< m1 >>
rect -7 5827 57 5897
<< viali >>
rect 0 5834 50 5890
<< locali >>
rect 2779 5827 2843 5897
<< m1 >>
rect 2779 5827 2843 5897
<< viali >>
rect 2786 5834 2836 5890
<< locali >>
rect 0 4170 2836 4226
<< locali >>
rect -7 4163 57 4233
<< m1 >>
rect -7 4163 57 4233
<< viali >>
rect 0 4170 50 4226
<< locali >>
rect 2779 4163 2843 4233
<< m1 >>
rect 2779 4163 2843 4233
<< viali >>
rect 2786 4170 2836 4226
<< labels >>
flabel m3 s 954 7913 984 8088 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m3 s 954 7113 984 7288 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 100 9840 2736 9890 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 0 9940 2836 9990 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m3 s 667 6713 697 7128 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
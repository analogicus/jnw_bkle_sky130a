magic
tech sky130A
magscale 1 1
timestamp 1748189726
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0  diff1_MP3<3> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 1940
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<2> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 1940
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<1> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 2340
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP3<0> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 2340
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<3> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 3140
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  diff1_MP4<3>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 3540
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP4<2> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 3140
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  diff1_MP4<2>_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 3540
box 0 0 576 240
use JNWATR_PCH_4C5F0  diff1_MP4<1> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 2740
box 0 0 576 400
use JNWATR_PCH_4C5F0  diff1_MP4<0> ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 2740
box 0 0 576 400
use JNWATR_PCH_4C5F0  mirror1_MP2 ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 1540
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  mirror1_MP2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 1300
box 0 0 576 240
use JNWATR_PCH_4C5F0  mirror1_MP1 ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 1540
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  mirror1_MP1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 1300
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN1 ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 440
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 840
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 3212 0 1 200
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN2 ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 440
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror2_MN2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 840
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mirror2_MN2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748189726
transform 1 0 2636 0 1 200
box 0 0 576 240
use JNWTR_RPPO16  bias1_RH1 ../JNW_TR_SKY130A
timestamp 1748189726
transform 1 0 200 0 1 200
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH2 ../JNW_TR_SKY130A
timestamp 1748189726
transform 1 0 200 0 1 3740
box 0 0 2236 1720
use JNWTR_RPPO16  bias1_RH3 ../JNW_TR_SKY130A
timestamp 1748189726
transform 1 0 200 0 1 1970
box 0 0 2236 1720
<< m2 >>
rect 3163 2123 3306 2153
<< m3 >>
rect 3163 2123 3193 2553
<< m2 >>
rect 3163 2523 3321 2553
<< m2 >>
rect 2715 2523 3321 2553
<< m2 >>
rect 2587 2523 2745 2553
<< m3 >>
rect 2587 2123 2617 2553
<< m2 >>
rect 2587 2123 2730 2153
<< m2 >>
rect 3156 2116 3200 2160
<< m3 >>
rect 3156 2116 3200 2160
<< via2 >>
rect 3163 2123 3193 2153
<< m2 >>
rect 3156 2516 3200 2560
<< m3 >>
rect 3156 2516 3200 2560
<< via2 >>
rect 3163 2523 3193 2553
<< m2 >>
rect 2580 2516 2624 2560
<< m3 >>
rect 2580 2516 2624 2560
<< via2 >>
rect 2587 2523 2617 2553
<< m2 >>
rect 2580 2116 2624 2160
<< m3 >>
rect 2580 2116 2624 2160
<< via2 >>
rect 2587 2123 2617 2153
<< m2 >>
rect 2587 3323 2730 3353
<< m3 >>
rect 2587 2923 2617 3353
<< m2 >>
rect 2587 2923 2745 2953
<< m2 >>
rect 2715 2923 3321 2953
<< m2 >>
rect 3163 2923 3321 2953
<< m3 >>
rect 3163 2923 3193 3353
<< m2 >>
rect 3163 3323 3306 3353
<< m2 >>
rect 2580 3316 2624 3360
<< m3 >>
rect 2580 3316 2624 3360
<< via2 >>
rect 2587 3323 2617 3353
<< m2 >>
rect 2580 2916 2624 2960
<< m3 >>
rect 2580 2916 2624 2960
<< via2 >>
rect 2587 2923 2617 2953
<< m2 >>
rect 3156 2916 3200 2960
<< m3 >>
rect 3156 2916 3200 2960
<< via2 >>
rect 3163 2923 3193 2953
<< m2 >>
rect 3156 3316 3200 3360
<< m3 >>
rect 3156 3316 3200 3360
<< via2 >>
rect 3163 3323 3193 3353
<< m2 >>
rect 2491 459 3018 489
<< m3 >>
rect 2491 459 2521 2793
<< m2 >>
rect 2491 2763 3033 2793
<< m3 >>
rect 3003 2763 3033 3193
<< m2 >>
rect 3003 3163 3609 3193
<< m3 >>
rect 3579 2778 3609 3193
<< m2 >>
rect 2484 452 2528 496
<< m3 >>
rect 2484 452 2528 496
<< via2 >>
rect 2491 459 2521 489
<< m2 >>
rect 2484 2756 2528 2800
<< m3 >>
rect 2484 2756 2528 2800
<< via2 >>
rect 2491 2763 2521 2793
<< m2 >>
rect 2996 2756 3040 2800
<< m3 >>
rect 2996 2756 3040 2800
<< via2 >>
rect 3003 2763 3033 2793
<< m2 >>
rect 2996 3156 3040 3200
<< m3 >>
rect 2996 3156 3040 3200
<< via2 >>
rect 3003 3163 3033 3193
<< m2 >>
rect 3572 3156 3616 3200
<< m3 >>
rect 3572 3156 3616 3200
<< via2 >>
rect 3579 3163 3609 3193
<< m2 >>
rect 2731 620 3322 650
<< m2 >>
rect 3164 620 3322 650
<< m3 >>
rect 3164 620 3194 1994
<< m2 >>
rect 3164 1964 3610 1994
<< m3 >>
rect 3580 1964 3610 2394
<< m2 >>
rect 3004 2364 3610 2394
<< m3 >>
rect 3004 1979 3034 2394
<< m2 >>
rect 3157 613 3201 657
<< m3 >>
rect 3157 613 3201 657
<< via2 >>
rect 3164 620 3194 650
<< m2 >>
rect 3157 1957 3201 2001
<< m3 >>
rect 3157 1957 3201 2001
<< via2 >>
rect 3164 1964 3194 1994
<< m2 >>
rect 3573 1957 3617 2001
<< m3 >>
rect 3573 1957 3617 2001
<< via2 >>
rect 3580 1964 3610 1994
<< m2 >>
rect 3573 2357 3617 2401
<< m3 >>
rect 3573 2357 3617 2401
<< via2 >>
rect 3580 2364 3610 2394
<< m2 >>
rect 2997 2357 3041 2401
<< m3 >>
rect 2997 2357 3041 2401
<< via2 >>
rect 3004 2364 3034 2394
<< m2 >>
rect 2396 1557 3019 1587
<< m3 >>
rect 2396 1557 2426 2275
<< m2 >>
rect 2396 2245 2842 2275
<< m2 >>
rect 2396 2245 2842 2275
<< m3 >>
rect 2396 2245 2426 2675
<< m2 >>
rect 2396 2645 2842 2675
<< m2 >>
rect 2396 2645 2842 2675
<< m3 >>
rect 2396 2645 2426 3075
<< m2 >>
rect 2396 3045 2842 3075
<< m2 >>
rect 2492 3045 2842 3075
<< m3 >>
rect 2492 3045 2522 3475
<< m2 >>
rect 2492 3445 2842 3475
<< m2 >>
rect 2812 3445 3418 3475
<< m2 >>
rect 3388 3445 3754 3475
<< m3 >>
rect 3724 3045 3754 3475
<< m2 >>
rect 3388 3045 3754 3075
<< m2 >>
rect 3388 3045 3754 3075
<< m3 >>
rect 3724 2645 3754 3075
<< m2 >>
rect 3388 2645 3754 2675
<< m2 >>
rect 3388 2645 3754 2675
<< m3 >>
rect 3724 2245 3754 2675
<< m2 >>
rect 3403 2245 3754 2275
<< m2 >>
rect 2389 1550 2433 1594
<< m3 >>
rect 2389 1550 2433 1594
<< via2 >>
rect 2396 1557 2426 1587
<< m2 >>
rect 2389 2238 2433 2282
<< m3 >>
rect 2389 2238 2433 2282
<< via2 >>
rect 2396 2245 2426 2275
<< m2 >>
rect 2389 2238 2433 2282
<< m3 >>
rect 2389 2238 2433 2282
<< via2 >>
rect 2396 2245 2426 2275
<< m2 >>
rect 2389 2638 2433 2682
<< m3 >>
rect 2389 2638 2433 2682
<< via2 >>
rect 2396 2645 2426 2675
<< m2 >>
rect 2389 2638 2433 2682
<< m3 >>
rect 2389 2638 2433 2682
<< via2 >>
rect 2396 2645 2426 2675
<< m2 >>
rect 2389 3038 2433 3082
<< m3 >>
rect 2389 3038 2433 3082
<< via2 >>
rect 2396 3045 2426 3075
<< m2 >>
rect 2485 3038 2529 3082
<< m3 >>
rect 2485 3038 2529 3082
<< via2 >>
rect 2492 3045 2522 3075
<< m2 >>
rect 2485 3438 2529 3482
<< m3 >>
rect 2485 3438 2529 3482
<< via2 >>
rect 2492 3445 2522 3475
<< m2 >>
rect 3717 3438 3761 3482
<< m3 >>
rect 3717 3438 3761 3482
<< via2 >>
rect 3724 3445 3754 3475
<< m2 >>
rect 3717 3038 3761 3082
<< m3 >>
rect 3717 3038 3761 3082
<< via2 >>
rect 3724 3045 3754 3075
<< m2 >>
rect 3717 3038 3761 3082
<< m3 >>
rect 3717 3038 3761 3082
<< via2 >>
rect 3724 3045 3754 3075
<< m2 >>
rect 3717 2638 3761 2682
<< m3 >>
rect 3717 2638 3761 2682
<< via2 >>
rect 3724 2645 3754 2675
<< m2 >>
rect 3717 2638 3761 2682
<< m3 >>
rect 3717 2638 3761 2682
<< via2 >>
rect 3724 2645 3754 2675
<< m2 >>
rect 3717 2238 3761 2282
<< m3 >>
rect 3717 2238 3761 2282
<< via2 >>
rect 3724 2245 3754 2275
<< m3 >>
rect 2170 1721 2200 1880
<< m2 >>
rect 2170 1850 2616 1880
<< m3 >>
rect 2586 1722 2616 1880
<< m2 >>
rect 2586 1722 2744 1752
<< m2 >>
rect 2714 1722 3305 1752
<< m2 >>
rect 2163 1843 2207 1887
<< m3 >>
rect 2163 1843 2207 1887
<< via2 >>
rect 2170 1850 2200 1880
<< m2 >>
rect 2579 1843 2623 1887
<< m3 >>
rect 2579 1843 2623 1887
<< via2 >>
rect 2586 1850 2616 1880
<< m2 >>
rect 2579 1715 2623 1759
<< m3 >>
rect 2579 1715 2623 1759
<< via2 >>
rect 2586 1722 2616 1752
<< m2 >>
rect 453 1703 2020 1733
<< m3 >>
rect 1990 1703 2020 5269
<< m2 >>
rect 1990 5239 2181 5269
<< m2 >>
rect 1983 1696 2027 1740
<< m3 >>
rect 1983 1696 2027 1740
<< via2 >>
rect 1990 1703 2020 1733
<< m2 >>
rect 1983 5232 2027 5276
<< m3 >>
rect 1983 5232 2027 5276
<< via2 >>
rect 1990 5239 2020 5269
<< m3 >>
rect 438 3689 468 5256
<< m2 >>
rect 438 3689 2196 3719
<< m3 >>
rect 2166 3480 2196 3719
<< m2 >>
rect 431 3682 475 3726
<< m3 >>
rect 431 3682 475 3726
<< via2 >>
rect 438 3689 468 3719
<< m2 >>
rect 2159 3682 2203 3726
<< m3 >>
rect 2159 3682 2203 3726
<< via2 >>
rect 2166 3689 2196 3719
<< locali >>
rect 100 5510 3980 5560
<< locali >>
rect 100 100 3980 150
<< m1 >>
rect 100 150 150 5510
<< m1 >>
rect 3930 150 3980 5510
<< locali >>
rect 93 5503 157 5567
<< m1 >>
rect 93 5503 157 5567
<< viali >>
rect 100 5510 150 5560
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 3923 5503 3987 5567
<< m1 >>
rect 3923 5503 3987 5567
<< viali >>
rect 3930 5510 3980 5560
<< locali >>
rect 3923 93 3987 157
<< m1 >>
rect 3923 93 3987 157
<< viali >>
rect 3930 100 3980 150
<< locali >>
rect 0 5610 4080 5660
<< locali >>
rect 0 0 4080 50
<< m1 >>
rect 0 50 50 5610
<< m1 >>
rect 4030 50 4080 5610
<< locali >>
rect -7 5603 57 5667
<< m1 >>
rect -7 5603 57 5667
<< viali >>
rect 0 5610 50 5660
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 4023 5603 4087 5667
<< m1 >>
rect 4023 5603 4087 5667
<< viali >>
rect 4030 5610 4080 5660
<< locali >>
rect 4023 -7 4087 57
<< m1 >>
rect 4023 -7 4087 57
<< viali >>
rect 4030 0 4080 50
<< locali >>
rect 208 3430 526 3550
<< locali >>
rect 100 1864 2436 1920
<< locali >>
rect 93 1857 157 1927
<< m1 >>
rect 93 1857 157 1927
<< viali >>
rect 100 1864 150 1920
<< locali >>
rect 100 200 2436 256
<< locali >>
rect 93 193 157 263
<< m1 >>
rect 93 193 157 263
<< viali >>
rect 100 200 150 256
<< locali >>
rect 100 5404 2436 5460
<< locali >>
rect 93 5397 157 5467
<< m1 >>
rect 93 5397 157 5467
<< viali >>
rect 100 5404 150 5460
<< locali >>
rect 100 3740 2436 3796
<< locali >>
rect 93 3733 157 3803
<< m1 >>
rect 93 3733 157 3803
<< viali >>
rect 100 3740 150 3796
<< locali >>
rect 100 3634 2436 3690
<< locali >>
rect 93 3627 157 3697
<< m1 >>
rect 93 3627 157 3697
<< viali >>
rect 100 3634 150 3690
<< locali >>
rect 100 1970 2436 2026
<< locali >>
rect 93 1963 157 2033
<< m1 >>
rect 93 1963 157 2033
<< viali >>
rect 100 1970 150 2026
<< locali >>
rect 2588 1840 2876 1880
<< locali >>
rect 3164 1840 3452 1880
<< locali >>
rect 3548 1720 3708 1760
<< locali >>
rect 3164 740 3452 780
<< locali >>
rect 3548 620 3708 660
<< locali >>
rect 2588 740 2876 780
<< locali >>
rect 2544 3612 4080 3708
<< locali >>
rect 4023 3605 4087 3715
<< m1 >>
rect 4023 3605 4087 3715
<< viali >>
rect 4030 3612 4080 3708
<< locali >>
rect 2544 1372 4080 1468
<< locali >>
rect 4023 1365 4087 1475
<< m1 >>
rect 4023 1365 4087 1475
<< viali >>
rect 4030 1372 4080 1468
<< locali >>
rect 2544 912 3980 1008
<< locali >>
rect 3923 905 3987 1015
<< m1 >>
rect 3923 905 3987 1015
<< viali >>
rect 3930 912 3980 1008
<< locali >>
rect 2544 272 3980 368
<< locali >>
rect 3923 265 3987 375
<< m1 >>
rect 3923 265 3987 375
<< viali >>
rect 3930 272 3980 368
<< m1 >>
rect 2709 2113 2755 2167
<< m2 >>
rect 2709 2113 2755 2167
<< via1 >>
rect 2716 2120 2748 2160
<< m1 >>
rect 3285 2113 3331 2167
<< m2 >>
rect 3285 2113 3331 2167
<< via1 >>
rect 3292 2120 3324 2160
<< m1 >>
rect 3285 2513 3331 2567
<< m2 >>
rect 3285 2513 3331 2567
<< via1 >>
rect 3292 2520 3324 2560
<< m1 >>
rect 3285 2513 3331 2567
<< m2 >>
rect 3285 2513 3331 2567
<< via1 >>
rect 3292 2520 3324 2560
<< m1 >>
rect 2709 2513 2755 2567
<< m2 >>
rect 2709 2513 2755 2567
<< via1 >>
rect 2716 2520 2748 2560
<< m1 >>
rect 2709 2513 2755 2567
<< m2 >>
rect 2709 2513 2755 2567
<< via1 >>
rect 2716 2520 2748 2560
<< m1 >>
rect 3285 3313 3331 3367
<< m2 >>
rect 3285 3313 3331 3367
<< via1 >>
rect 3292 3320 3324 3360
<< m1 >>
rect 2709 3313 2755 3367
<< m2 >>
rect 2709 3313 2755 3367
<< via1 >>
rect 2716 3320 2748 3360
<< m1 >>
rect 3285 2913 3331 2967
<< m2 >>
rect 3285 2913 3331 2967
<< via1 >>
rect 3292 2920 3324 2960
<< m1 >>
rect 3285 2913 3331 2967
<< m2 >>
rect 3285 2913 3331 2967
<< via1 >>
rect 3292 2920 3324 2960
<< m1 >>
rect 2709 2913 2755 2967
<< m2 >>
rect 2709 2913 2755 2967
<< via1 >>
rect 2716 2920 2748 2960
<< m1 >>
rect 2709 2913 2755 2967
<< m2 >>
rect 2709 2913 2755 2967
<< via1 >>
rect 2716 2920 2748 2960
<< m1 >>
rect 3541 3153 3651 3207
<< m2 >>
rect 3541 3153 3651 3207
<< via1 >>
rect 3548 3160 3644 3200
<< m1 >>
rect 3541 3153 3651 3207
<< m2 >>
rect 3541 3153 3651 3207
<< m3 >>
rect 3541 3153 3651 3207
<< via2 >>
rect 3548 3160 3644 3200
<< via1 >>
rect 3548 3160 3644 3200
<< m1 >>
rect 2965 3153 3075 3207
<< m2 >>
rect 2965 3153 3075 3207
<< m3 >>
rect 2965 3153 3075 3207
<< via2 >>
rect 2972 3160 3068 3200
<< via1 >>
rect 2972 3160 3068 3200
<< m1 >>
rect 2965 3153 3075 3207
<< m2 >>
rect 2965 3153 3075 3207
<< via1 >>
rect 2972 3160 3068 3200
<< m1 >>
rect 3541 2753 3651 2807
<< m2 >>
rect 3541 2753 3651 2807
<< m3 >>
rect 3541 2753 3651 2807
<< via2 >>
rect 3548 2760 3644 2800
<< via1 >>
rect 3548 2760 3644 2800
<< m1 >>
rect 2965 2753 3075 2807
<< m2 >>
rect 2965 2753 3075 2807
<< via1 >>
rect 2972 2760 3068 2800
<< m1 >>
rect 2965 2753 3075 2807
<< m2 >>
rect 2965 2753 3075 2807
<< m3 >>
rect 2965 2753 3075 2807
<< via2 >>
rect 2972 2760 3068 2800
<< via1 >>
rect 2972 2760 3068 2800
<< m1 >>
rect 2965 453 3075 507
<< m2 >>
rect 2965 453 3075 507
<< via1 >>
rect 2972 460 3068 500
<< m1 >>
rect 2965 1953 3075 2007
<< m2 >>
rect 2965 1953 3075 2007
<< m3 >>
rect 2965 1953 3075 2007
<< via2 >>
rect 2972 1960 3068 2000
<< via1 >>
rect 2972 1960 3068 2000
<< m1 >>
rect 3541 1953 3651 2007
<< m2 >>
rect 3541 1953 3651 2007
<< via1 >>
rect 3548 1960 3644 2000
<< m1 >>
rect 3541 1953 3651 2007
<< m2 >>
rect 3541 1953 3651 2007
<< m3 >>
rect 3541 1953 3651 2007
<< via2 >>
rect 3548 1960 3644 2000
<< via1 >>
rect 3548 1960 3644 2000
<< m1 >>
rect 3541 2353 3651 2407
<< m2 >>
rect 3541 2353 3651 2407
<< m3 >>
rect 3541 2353 3651 2407
<< via2 >>
rect 3548 2360 3644 2400
<< via1 >>
rect 3548 2360 3644 2400
<< m1 >>
rect 3541 2353 3651 2407
<< m2 >>
rect 3541 2353 3651 2407
<< via1 >>
rect 3548 2360 3644 2400
<< m1 >>
rect 2965 2353 3075 2407
<< m2 >>
rect 2965 2353 3075 2407
<< via1 >>
rect 2972 2360 3068 2400
<< m1 >>
rect 2965 2353 3075 2407
<< m2 >>
rect 2965 2353 3075 2407
<< m3 >>
rect 2965 2353 3075 2407
<< via2 >>
rect 2972 2360 3068 2400
<< via1 >>
rect 2972 2360 3068 2400
<< m1 >>
rect 3285 613 3331 667
<< m2 >>
rect 3285 613 3331 667
<< via1 >>
rect 3292 620 3324 660
<< m1 >>
rect 3285 613 3331 667
<< m2 >>
rect 3285 613 3331 667
<< via1 >>
rect 3292 620 3324 660
<< m1 >>
rect 2709 613 2755 667
<< m2 >>
rect 2709 613 2755 667
<< via1 >>
rect 2716 620 2748 660
<< m1 >>
rect 2773 2233 2883 2287
<< m2 >>
rect 2773 2233 2883 2287
<< via1 >>
rect 2780 2240 2876 2280
<< m1 >>
rect 2773 2233 2883 2287
<< m2 >>
rect 2773 2233 2883 2287
<< via1 >>
rect 2780 2240 2876 2280
<< m1 >>
rect 3349 2233 3459 2287
<< m2 >>
rect 3349 2233 3459 2287
<< via1 >>
rect 3356 2240 3452 2280
<< m1 >>
rect 3349 2633 3459 2687
<< m2 >>
rect 3349 2633 3459 2687
<< via1 >>
rect 3356 2640 3452 2680
<< m1 >>
rect 3349 2633 3459 2687
<< m2 >>
rect 3349 2633 3459 2687
<< via1 >>
rect 3356 2640 3452 2680
<< m1 >>
rect 2773 2633 2883 2687
<< m2 >>
rect 2773 2633 2883 2687
<< via1 >>
rect 2780 2640 2876 2680
<< m1 >>
rect 2773 2633 2883 2687
<< m2 >>
rect 2773 2633 2883 2687
<< via1 >>
rect 2780 2640 2876 2680
<< m1 >>
rect 3349 3433 3459 3487
<< m2 >>
rect 3349 3433 3459 3487
<< via1 >>
rect 3356 3440 3452 3480
<< m1 >>
rect 3349 3433 3459 3487
<< m2 >>
rect 3349 3433 3459 3487
<< via1 >>
rect 3356 3440 3452 3480
<< m1 >>
rect 2773 3433 2883 3487
<< m2 >>
rect 2773 3433 2883 3487
<< via1 >>
rect 2780 3440 2876 3480
<< m1 >>
rect 2773 3433 2883 3487
<< m2 >>
rect 2773 3433 2883 3487
<< via1 >>
rect 2780 3440 2876 3480
<< m1 >>
rect 3349 3033 3459 3087
<< m2 >>
rect 3349 3033 3459 3087
<< via1 >>
rect 3356 3040 3452 3080
<< m1 >>
rect 3349 3033 3459 3087
<< m2 >>
rect 3349 3033 3459 3087
<< via1 >>
rect 3356 3040 3452 3080
<< m1 >>
rect 2773 3033 2883 3087
<< m2 >>
rect 2773 3033 2883 3087
<< via1 >>
rect 2780 3040 2876 3080
<< m1 >>
rect 2773 3033 2883 3087
<< m2 >>
rect 2773 3033 2883 3087
<< via1 >>
rect 2780 3040 2876 3080
<< m1 >>
rect 2965 1553 3075 1607
<< m2 >>
rect 2965 1553 3075 1607
<< via1 >>
rect 2972 1560 3068 1600
<< m1 >>
rect 2709 1713 2755 1767
<< m2 >>
rect 2709 1713 2755 1767
<< via1 >>
rect 2716 1720 2748 1760
<< m1 >>
rect 2709 1713 2755 1767
<< m2 >>
rect 2709 1713 2755 1767
<< via1 >>
rect 2716 1720 2748 1760
<< m1 >>
rect 3285 1713 3331 1767
<< m2 >>
rect 3285 1713 3331 1767
<< via1 >>
rect 3292 1720 3324 1760
<< locali >>
rect 2103 1653 2261 1787
<< m1 >>
rect 2103 1653 2261 1787
<< m2 >>
rect 2103 1653 2261 1787
<< m3 >>
rect 2103 1653 2261 1787
<< via2 >>
rect 2110 1660 2254 1780
<< via1 >>
rect 2110 1660 2254 1780
<< viali >>
rect 2110 1660 2254 1780
<< locali >>
rect 375 1653 533 1787
<< m1 >>
rect 375 1653 533 1787
<< m2 >>
rect 375 1653 533 1787
<< via1 >>
rect 382 1660 526 1780
<< viali >>
rect 382 1660 526 1780
<< locali >>
rect 2103 5193 2261 5327
<< m1 >>
rect 2103 5193 2261 5327
<< m2 >>
rect 2103 5193 2261 5327
<< via1 >>
rect 2110 5200 2254 5320
<< viali >>
rect 2110 5200 2254 5320
<< locali >>
rect 375 5193 533 5327
<< m1 >>
rect 375 5193 533 5327
<< m2 >>
rect 375 5193 533 5327
<< m3 >>
rect 375 5193 533 5327
<< via2 >>
rect 382 5200 526 5320
<< via1 >>
rect 382 5200 526 5320
<< viali >>
rect 382 5200 526 5320
<< locali >>
rect 2103 3423 2261 3557
<< m1 >>
rect 2103 3423 2261 3557
<< m2 >>
rect 2103 3423 2261 3557
<< m3 >>
rect 2103 3423 2261 3557
<< via2 >>
rect 2110 3430 2254 3550
<< via1 >>
rect 2110 3430 2254 3550
<< viali >>
rect 2110 3430 2254 3550
<< labels >>
flabel m2 s 3163 2123 3306 2153 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 2587 3323 2730 3353 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 0 5610 4080 5660 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 100 5510 3980 5560 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m2 s 2491 459 3018 489 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
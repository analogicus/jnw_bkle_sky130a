magic
tech sky130A
magscale 1 1
timestamp 1748755918
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0  df1_MP3<3> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 1540
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  df1_MP3<3>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 1300
box 0 0 576 240
use JNWATR_PCH_4C5F0  df1_MP3<2> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 1540
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  df1_MP3<2>_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 1300
box 0 0 576 240
use JNWATR_PCH_4C5F0  df1_MP3<1> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 1940
box 0 0 576 400
use JNWATR_PCH_4C5F0  df1_MP3<0> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 1940
box 0 0 576 400
use JNWATR_PCH_4C5F0  df1_MP4<3> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 2340
box 0 0 576 400
use JNWATR_PCH_4C5F0  df1_MP4<2> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 2340
box 0 0 576 400
use JNWATR_PCH_4C5F0  df1_MP4<1> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 2740
box 0 0 576 400
use JNWATR_PCH_4C5F0  df1_MP4<0> ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 2740
box 0 0 576 400
use JNWATR_PCH_4C5F0  mr1_MP2 ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 3140
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mr1_MP2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 3540
box 0 0 576 240
use JNWATR_PCH_4C5F0  mr1_MP1 ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 3140
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  mr1_MP1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 3540
box 0 0 576 240
use JNWATR_NCH_4C5F0  mr2_MN1 ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 440
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mr2_MN1_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 840
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mr2_MN1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 3212 0 1 200
box 0 0 576 240
use JNWATR_NCH_4C5F0  mr2_MN2 ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 440
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mr2_MN2_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 840
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT  mr2_MN2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748755918
transform 1 0 2636 0 1 200
box 0 0 576 240
use JNWTR_RPPO16  bs1_RH1 ../JNW_TR_SKY130A
timestamp 1748755918
transform 1 0 200 0 1 200
box 0 0 2236 1720
use JNWTR_RPPO16  bs1_RH2 ../JNW_TR_SKY130A
timestamp 1748755918
transform 1 0 200 0 1 3740
box 0 0 2236 1720
use JNWTR_RPPO16  bs1_RH3 ../JNW_TR_SKY130A
timestamp 1748755918
transform 1 0 200 0 1 1970
box 0 0 2236 1720
<< m2 >>
rect 3163 1723 3306 1753
<< m3 >>
rect 3163 1723 3193 2153
<< m2 >>
rect 3163 2123 3321 2153
<< m2 >>
rect 2715 2123 3321 2153
<< m2 >>
rect 2587 2123 2745 2153
<< m3 >>
rect 2587 1723 2617 2153
<< m2 >>
rect 2587 1723 2730 1753
<< m2 >>
rect 3156 1716 3200 1760
<< m3 >>
rect 3156 1716 3200 1760
<< via2 >>
rect 3163 1723 3193 1753
<< m2 >>
rect 3156 2116 3200 2160
<< m3 >>
rect 3156 2116 3200 2160
<< via2 >>
rect 3163 2123 3193 2153
<< m2 >>
rect 2580 2116 2624 2160
<< m3 >>
rect 2580 2116 2624 2160
<< via2 >>
rect 2587 2123 2617 2153
<< m2 >>
rect 2580 1716 2624 1760
<< m3 >>
rect 2580 1716 2624 1760
<< via2 >>
rect 2587 1723 2617 1753
<< m2 >>
rect 3163 2523 3306 2553
<< m3 >>
rect 3163 2523 3193 2953
<< m2 >>
rect 3163 2923 3321 2953
<< m2 >>
rect 2715 2923 3321 2953
<< m2 >>
rect 2587 2923 2745 2953
<< m3 >>
rect 2587 2523 2617 2953
<< m2 >>
rect 2587 2523 2730 2553
<< m2 >>
rect 3156 2516 3200 2560
<< m3 >>
rect 3156 2516 3200 2560
<< via2 >>
rect 3163 2523 3193 2553
<< m2 >>
rect 3156 2916 3200 2960
<< m3 >>
rect 3156 2916 3200 2960
<< via2 >>
rect 3163 2923 3193 2953
<< m2 >>
rect 2580 2916 2624 2960
<< m3 >>
rect 2580 2916 2624 2960
<< via2 >>
rect 2587 2923 2617 2953
<< m2 >>
rect 2580 2516 2624 2560
<< m3 >>
rect 2580 2516 2624 2560
<< via2 >>
rect 2587 2523 2617 2553
<< m2 >>
rect 2491 459 3018 489
<< m3 >>
rect 2491 459 2521 2393
<< m2 >>
rect 2491 2363 3033 2393
<< m3 >>
rect 3003 2363 3033 2793
<< m2 >>
rect 3003 2763 3609 2793
<< m3 >>
rect 3579 2378 3609 2793
<< m2 >>
rect 2484 452 2528 496
<< m3 >>
rect 2484 452 2528 496
<< via2 >>
rect 2491 459 2521 489
<< m2 >>
rect 2484 2356 2528 2400
<< m3 >>
rect 2484 2356 2528 2400
<< via2 >>
rect 2491 2363 2521 2393
<< m2 >>
rect 2996 2356 3040 2400
<< m3 >>
rect 2996 2356 3040 2400
<< via2 >>
rect 3003 2363 3033 2393
<< m2 >>
rect 2996 2756 3040 2800
<< m3 >>
rect 2996 2756 3040 2800
<< via2 >>
rect 3003 2763 3033 2793
<< m2 >>
rect 3572 2756 3616 2800
<< m3 >>
rect 3572 2756 3616 2800
<< via2 >>
rect 3579 2763 3609 2793
<< m2 >>
rect 2731 620 3322 650
<< m2 >>
rect 3292 620 3610 650
<< m3 >>
rect 3580 620 3610 1594
<< m3 >>
rect 3580 1564 3610 1994
<< m2 >>
rect 3004 1964 3610 1994
<< m3 >>
rect 3004 1579 3034 1994
<< m2 >>
rect 3573 613 3617 657
<< m3 >>
rect 3573 613 3617 657
<< via2 >>
rect 3580 620 3610 650
<< m2 >>
rect 3573 1957 3617 2001
<< m3 >>
rect 3573 1957 3617 2001
<< via2 >>
rect 3580 1964 3610 1994
<< m2 >>
rect 2997 1957 3041 2001
<< m3 >>
rect 2997 1957 3041 2001
<< via2 >>
rect 3004 1964 3034 1994
<< m2 >>
rect 2844 3157 3019 3187
<< m3 >>
rect 2844 2773 2874 3187
<< m2 >>
rect 2684 2773 2874 2803
<< m3 >>
rect 2684 2645 2714 2803
<< m2 >>
rect 2684 2645 2842 2675
<< m2 >>
rect 2860 3045 3418 3075
<< m2 >>
rect 3388 3045 3754 3075
<< m3 >>
rect 3724 2645 3754 3075
<< m2 >>
rect 3388 2645 3754 2675
<< m2 >>
rect 3388 2645 3754 2675
<< m3 >>
rect 3724 2245 3754 2675
<< m2 >>
rect 3388 2245 3754 2275
<< m2 >>
rect 3388 2245 3754 2275
<< m3 >>
rect 3724 1845 3754 2275
<< m2 >>
rect 3388 1845 3754 1875
<< m2 >>
rect 2812 1845 3418 1875
<< m2 >>
rect 2396 1845 2842 1875
<< m3 >>
rect 2396 1845 2426 2275
<< m2 >>
rect 2396 2245 2827 2275
<< m2 >>
rect 2837 3150 2881 3194
<< m3 >>
rect 2837 3150 2881 3194
<< via2 >>
rect 2844 3157 2874 3187
<< m2 >>
rect 2837 2766 2881 2810
<< m3 >>
rect 2837 2766 2881 2810
<< via2 >>
rect 2844 2773 2874 2803
<< m2 >>
rect 2677 2766 2721 2810
<< m3 >>
rect 2677 2766 2721 2810
<< via2 >>
rect 2684 2773 2714 2803
<< m2 >>
rect 2677 2638 2721 2682
<< m3 >>
rect 2677 2638 2721 2682
<< via2 >>
rect 2684 2645 2714 2675
<< m2 >>
rect 3717 3038 3761 3082
<< m3 >>
rect 3717 3038 3761 3082
<< via2 >>
rect 3724 3045 3754 3075
<< m2 >>
rect 3717 2638 3761 2682
<< m3 >>
rect 3717 2638 3761 2682
<< via2 >>
rect 3724 2645 3754 2675
<< m2 >>
rect 3717 2638 3761 2682
<< m3 >>
rect 3717 2638 3761 2682
<< via2 >>
rect 3724 2645 3754 2675
<< m2 >>
rect 3717 2238 3761 2282
<< m3 >>
rect 3717 2238 3761 2282
<< via2 >>
rect 3724 2245 3754 2275
<< m2 >>
rect 3717 2238 3761 2282
<< m3 >>
rect 3717 2238 3761 2282
<< via2 >>
rect 3724 2245 3754 2275
<< m2 >>
rect 3717 1838 3761 1882
<< m3 >>
rect 3717 1838 3761 1882
<< via2 >>
rect 3724 1845 3754 1875
<< m2 >>
rect 2389 1838 2433 1882
<< m3 >>
rect 2389 1838 2433 1882
<< via2 >>
rect 2396 1845 2426 1875
<< m2 >>
rect 2389 2238 2433 2282
<< m3 >>
rect 2389 2238 2433 2282
<< via2 >>
rect 2396 2245 2426 2275
<< m3 >>
rect 2170 1721 2200 3176
<< m2 >>
rect 2170 3146 2392 3176
<< m3 >>
rect 2362 3146 2392 3352
<< m2 >>
rect 2362 3322 2744 3352
<< m2 >>
rect 2714 3322 3305 3352
<< m2 >>
rect 2163 3139 2207 3183
<< m3 >>
rect 2163 3139 2207 3183
<< via2 >>
rect 2170 3146 2200 3176
<< m2 >>
rect 2355 3139 2399 3183
<< m3 >>
rect 2355 3139 2399 3183
<< via2 >>
rect 2362 3146 2392 3176
<< m2 >>
rect 2355 3315 2399 3359
<< m3 >>
rect 2355 3315 2399 3359
<< via2 >>
rect 2362 3322 2392 3352
<< m2 >>
rect 453 1703 2020 1733
<< m3 >>
rect 1990 1703 2020 5269
<< m2 >>
rect 1990 5239 2181 5269
<< m2 >>
rect 1983 1696 2027 1740
<< m3 >>
rect 1983 1696 2027 1740
<< via2 >>
rect 1990 1703 2020 1733
<< m2 >>
rect 1983 5232 2027 5276
<< m3 >>
rect 1983 5232 2027 5276
<< via2 >>
rect 1990 5239 2020 5269
<< m3 >>
rect 438 3689 468 5256
<< m2 >>
rect 438 3689 2196 3719
<< m3 >>
rect 2166 3480 2196 3719
<< m2 >>
rect 431 3682 475 3726
<< m3 >>
rect 431 3682 475 3726
<< via2 >>
rect 438 3689 468 3719
<< m2 >>
rect 2159 3682 2203 3726
<< m3 >>
rect 2159 3682 2203 3726
<< via2 >>
rect 2166 3689 2196 3719
<< locali >>
rect 100 5510 3980 5560
<< locali >>
rect 100 100 3980 150
<< m1 >>
rect 100 150 150 5510
<< m1 >>
rect 3930 150 3980 5510
<< locali >>
rect 93 5503 157 5567
<< m1 >>
rect 93 5503 157 5567
<< viali >>
rect 100 5510 150 5560
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 3923 5503 3987 5567
<< m1 >>
rect 3923 5503 3987 5567
<< viali >>
rect 3930 5510 3980 5560
<< locali >>
rect 3923 93 3987 157
<< m1 >>
rect 3923 93 3987 157
<< viali >>
rect 3930 100 3980 150
<< locali >>
rect 0 5610 4080 5660
<< locali >>
rect 0 0 4080 50
<< m1 >>
rect 0 50 50 5610
<< m1 >>
rect 4030 50 4080 5610
<< locali >>
rect -7 5603 57 5667
<< m1 >>
rect -7 5603 57 5667
<< viali >>
rect 0 5610 50 5660
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 4023 5603 4087 5667
<< m1 >>
rect 4023 5603 4087 5667
<< viali >>
rect 4030 5610 4080 5660
<< locali >>
rect 4023 -7 4087 57
<< m1 >>
rect 4023 -7 4087 57
<< viali >>
rect 4030 0 4080 50
<< locali >>
rect 208 3430 526 3550
<< locali >>
rect 100 1864 2436 1920
<< locali >>
rect 93 1857 157 1927
<< m1 >>
rect 93 1857 157 1927
<< viali >>
rect 100 1864 150 1920
<< locali >>
rect 100 200 2436 256
<< locali >>
rect 93 193 157 263
<< m1 >>
rect 93 193 157 263
<< viali >>
rect 100 200 150 256
<< locali >>
rect 100 5404 2436 5460
<< locali >>
rect 93 5397 157 5467
<< m1 >>
rect 93 5397 157 5467
<< viali >>
rect 100 5404 150 5460
<< locali >>
rect 100 3740 2436 3796
<< locali >>
rect 93 3733 157 3803
<< m1 >>
rect 93 3733 157 3803
<< viali >>
rect 100 3740 150 3796
<< locali >>
rect 100 3634 2436 3690
<< locali >>
rect 93 3627 157 3697
<< m1 >>
rect 93 3627 157 3697
<< viali >>
rect 100 3634 150 3690
<< locali >>
rect 100 1970 2436 2026
<< locali >>
rect 93 1963 157 2033
<< m1 >>
rect 93 1963 157 2033
<< viali >>
rect 100 1970 150 2026
<< locali >>
rect 2588 3440 2876 3480
<< locali >>
rect 3164 3440 3452 3480
<< locali >>
rect 3548 3320 3708 3360
<< locali >>
rect 3164 740 3452 780
<< locali >>
rect 3548 620 3708 660
<< locali >>
rect 2588 740 2876 780
<< locali >>
rect 2544 1372 4080 1468
<< locali >>
rect 4023 1365 4087 1475
<< m1 >>
rect 4023 1365 4087 1475
<< viali >>
rect 4030 1372 4080 1468
<< locali >>
rect 2544 3612 4080 3708
<< locali >>
rect 4023 3605 4087 3715
<< m1 >>
rect 4023 3605 4087 3715
<< viali >>
rect 4030 3612 4080 3708
<< locali >>
rect 2544 912 3980 1008
<< locali >>
rect 3923 905 3987 1015
<< m1 >>
rect 3923 905 3987 1015
<< viali >>
rect 3930 912 3980 1008
<< locali >>
rect 2544 272 3980 368
<< locali >>
rect 3923 265 3987 375
<< m1 >>
rect 3923 265 3987 375
<< viali >>
rect 3930 272 3980 368
<< m1 >>
rect 2709 1713 2755 1767
<< m2 >>
rect 2709 1713 2755 1767
<< via1 >>
rect 2716 1720 2748 1760
<< m1 >>
rect 3285 1713 3331 1767
<< m2 >>
rect 3285 1713 3331 1767
<< via1 >>
rect 3292 1720 3324 1760
<< m1 >>
rect 3285 2113 3331 2167
<< m2 >>
rect 3285 2113 3331 2167
<< via1 >>
rect 3292 2120 3324 2160
<< m1 >>
rect 3285 2113 3331 2167
<< m2 >>
rect 3285 2113 3331 2167
<< via1 >>
rect 3292 2120 3324 2160
<< m1 >>
rect 2709 2113 2755 2167
<< m2 >>
rect 2709 2113 2755 2167
<< via1 >>
rect 2716 2120 2748 2160
<< m1 >>
rect 2709 2113 2755 2167
<< m2 >>
rect 2709 2113 2755 2167
<< via1 >>
rect 2716 2120 2748 2160
<< m1 >>
rect 2709 2513 2755 2567
<< m2 >>
rect 2709 2513 2755 2567
<< via1 >>
rect 2716 2520 2748 2560
<< m1 >>
rect 3285 2513 3331 2567
<< m2 >>
rect 3285 2513 3331 2567
<< via1 >>
rect 3292 2520 3324 2560
<< m1 >>
rect 2709 2913 2755 2967
<< m2 >>
rect 2709 2913 2755 2967
<< via1 >>
rect 2716 2920 2748 2960
<< m1 >>
rect 2709 2913 2755 2967
<< m2 >>
rect 2709 2913 2755 2967
<< via1 >>
rect 2716 2920 2748 2960
<< m1 >>
rect 3285 2913 3331 2967
<< m2 >>
rect 3285 2913 3331 2967
<< via1 >>
rect 3292 2920 3324 2960
<< m1 >>
rect 3285 2913 3331 2967
<< m2 >>
rect 3285 2913 3331 2967
<< via1 >>
rect 3292 2920 3324 2960
<< m1 >>
rect 2965 2353 3075 2407
<< m2 >>
rect 2965 2353 3075 2407
<< via1 >>
rect 2972 2360 3068 2400
<< m1 >>
rect 2965 2353 3075 2407
<< m2 >>
rect 2965 2353 3075 2407
<< m3 >>
rect 2965 2353 3075 2407
<< via2 >>
rect 2972 2360 3068 2400
<< via1 >>
rect 2972 2360 3068 2400
<< m1 >>
rect 3541 2353 3651 2407
<< m2 >>
rect 3541 2353 3651 2407
<< m3 >>
rect 3541 2353 3651 2407
<< via2 >>
rect 3548 2360 3644 2400
<< via1 >>
rect 3548 2360 3644 2400
<< m1 >>
rect 2965 2753 3075 2807
<< m2 >>
rect 2965 2753 3075 2807
<< m3 >>
rect 2965 2753 3075 2807
<< via2 >>
rect 2972 2760 3068 2800
<< via1 >>
rect 2972 2760 3068 2800
<< m1 >>
rect 2965 2753 3075 2807
<< m2 >>
rect 2965 2753 3075 2807
<< via1 >>
rect 2972 2760 3068 2800
<< m1 >>
rect 3541 2753 3651 2807
<< m2 >>
rect 3541 2753 3651 2807
<< via1 >>
rect 3548 2760 3644 2800
<< m1 >>
rect 3541 2753 3651 2807
<< m2 >>
rect 3541 2753 3651 2807
<< m3 >>
rect 3541 2753 3651 2807
<< via2 >>
rect 3548 2760 3644 2800
<< via1 >>
rect 3548 2760 3644 2800
<< m1 >>
rect 2965 453 3075 507
<< m2 >>
rect 2965 453 3075 507
<< via1 >>
rect 2972 460 3068 500
<< m1 >>
rect 2965 1553 3075 1607
<< m2 >>
rect 2965 1553 3075 1607
<< m3 >>
rect 2965 1553 3075 1607
<< via2 >>
rect 2972 1560 3068 1600
<< via1 >>
rect 2972 1560 3068 1600
<< m1 >>
rect 3541 1553 3651 1607
<< m2 >>
rect 3541 1553 3651 1607
<< m3 >>
rect 3541 1553 3651 1607
<< via2 >>
rect 3548 1560 3644 1600
<< via1 >>
rect 3548 1560 3644 1600
<< m1 >>
rect 3541 1553 3651 1607
<< m2 >>
rect 3541 1553 3651 1607
<< m3 >>
rect 3541 1553 3651 1607
<< via2 >>
rect 3548 1560 3644 1600
<< via1 >>
rect 3548 1560 3644 1600
<< m1 >>
rect 3541 1953 3651 2007
<< m2 >>
rect 3541 1953 3651 2007
<< m3 >>
rect 3541 1953 3651 2007
<< via2 >>
rect 3548 1960 3644 2000
<< via1 >>
rect 3548 1960 3644 2000
<< m1 >>
rect 3541 1953 3651 2007
<< m2 >>
rect 3541 1953 3651 2007
<< via1 >>
rect 3548 1960 3644 2000
<< m1 >>
rect 2965 1953 3075 2007
<< m2 >>
rect 2965 1953 3075 2007
<< via1 >>
rect 2972 1960 3068 2000
<< m1 >>
rect 2965 1953 3075 2007
<< m2 >>
rect 2965 1953 3075 2007
<< m3 >>
rect 2965 1953 3075 2007
<< via2 >>
rect 2972 1960 3068 2000
<< via1 >>
rect 2972 1960 3068 2000
<< m1 >>
rect 3285 613 3331 667
<< m2 >>
rect 3285 613 3331 667
<< via1 >>
rect 3292 620 3324 660
<< m1 >>
rect 3285 613 3331 667
<< m2 >>
rect 3285 613 3331 667
<< via1 >>
rect 3292 620 3324 660
<< m1 >>
rect 2709 613 2755 667
<< m2 >>
rect 2709 613 2755 667
<< via1 >>
rect 2716 620 2748 660
<< m1 >>
rect 2773 1833 2883 1887
<< m2 >>
rect 2773 1833 2883 1887
<< via1 >>
rect 2780 1840 2876 1880
<< m1 >>
rect 2773 1833 2883 1887
<< m2 >>
rect 2773 1833 2883 1887
<< via1 >>
rect 2780 1840 2876 1880
<< m1 >>
rect 3349 1833 3459 1887
<< m2 >>
rect 3349 1833 3459 1887
<< via1 >>
rect 3356 1840 3452 1880
<< m1 >>
rect 3349 1833 3459 1887
<< m2 >>
rect 3349 1833 3459 1887
<< via1 >>
rect 3356 1840 3452 1880
<< m1 >>
rect 3349 2233 3459 2287
<< m2 >>
rect 3349 2233 3459 2287
<< via1 >>
rect 3356 2240 3452 2280
<< m1 >>
rect 3349 2233 3459 2287
<< m2 >>
rect 3349 2233 3459 2287
<< via1 >>
rect 3356 2240 3452 2280
<< m1 >>
rect 2773 2233 2883 2287
<< m2 >>
rect 2773 2233 2883 2287
<< via1 >>
rect 2780 2240 2876 2280
<< m1 >>
rect 2773 2633 2883 2687
<< m2 >>
rect 2773 2633 2883 2687
<< via1 >>
rect 2780 2640 2876 2680
<< m1 >>
rect 3349 2633 3459 2687
<< m2 >>
rect 3349 2633 3459 2687
<< via1 >>
rect 3356 2640 3452 2680
<< m1 >>
rect 3349 2633 3459 2687
<< m2 >>
rect 3349 2633 3459 2687
<< via1 >>
rect 3356 2640 3452 2680
<< m1 >>
rect 2773 3033 2883 3087
<< m2 >>
rect 2773 3033 2883 3087
<< m3 >>
rect 2773 3033 2883 3087
<< via2 >>
rect 2780 3040 2876 3080
<< via1 >>
rect 2780 3040 2876 3080
<< m1 >>
rect 2773 3033 2883 3087
<< m2 >>
rect 2773 3033 2883 3087
<< via1 >>
rect 2780 3040 2876 3080
<< m1 >>
rect 3349 3033 3459 3087
<< m2 >>
rect 3349 3033 3459 3087
<< via1 >>
rect 3356 3040 3452 3080
<< m1 >>
rect 3349 3033 3459 3087
<< m2 >>
rect 3349 3033 3459 3087
<< via1 >>
rect 3356 3040 3452 3080
<< m1 >>
rect 2965 3153 3075 3207
<< m2 >>
rect 2965 3153 3075 3207
<< via1 >>
rect 2972 3160 3068 3200
<< m1 >>
rect 2709 3313 2755 3367
<< m2 >>
rect 2709 3313 2755 3367
<< via1 >>
rect 2716 3320 2748 3360
<< m1 >>
rect 2709 3313 2755 3367
<< m2 >>
rect 2709 3313 2755 3367
<< via1 >>
rect 2716 3320 2748 3360
<< m1 >>
rect 3285 3313 3331 3367
<< m2 >>
rect 3285 3313 3331 3367
<< via1 >>
rect 3292 3320 3324 3360
<< locali >>
rect 2103 1653 2261 1787
<< m1 >>
rect 2103 1653 2261 1787
<< m2 >>
rect 2103 1653 2261 1787
<< m3 >>
rect 2103 1653 2261 1787
<< via2 >>
rect 2110 1660 2254 1780
<< via1 >>
rect 2110 1660 2254 1780
<< viali >>
rect 2110 1660 2254 1780
<< locali >>
rect 375 1653 533 1787
<< m1 >>
rect 375 1653 533 1787
<< m2 >>
rect 375 1653 533 1787
<< via1 >>
rect 382 1660 526 1780
<< viali >>
rect 382 1660 526 1780
<< locali >>
rect 2103 5193 2261 5327
<< m1 >>
rect 2103 5193 2261 5327
<< m2 >>
rect 2103 5193 2261 5327
<< via1 >>
rect 2110 5200 2254 5320
<< viali >>
rect 2110 5200 2254 5320
<< locali >>
rect 375 5193 533 5327
<< m1 >>
rect 375 5193 533 5327
<< m2 >>
rect 375 5193 533 5327
<< m3 >>
rect 375 5193 533 5327
<< via2 >>
rect 382 5200 526 5320
<< via1 >>
rect 382 5200 526 5320
<< viali >>
rect 382 5200 526 5320
<< locali >>
rect 2103 3423 2261 3557
<< m1 >>
rect 2103 3423 2261 3557
<< m2 >>
rect 2103 3423 2261 3557
<< m3 >>
rect 2103 3423 2261 3557
<< via2 >>
rect 2110 3430 2254 3550
<< via1 >>
rect 2110 3430 2254 3550
<< viali >>
rect 2110 3430 2254 3550
<< labels >>
flabel m2 s 3163 1723 3306 1753 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 3163 2523 3306 2553 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 0 5610 4080 5660 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 100 5510 3980 5560 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m2 s 2491 459 3018 489 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1743432408
<< checkpaint >>
rect 0 0 0 0
use JNWATR_PCH_4C1F2 diff1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 1600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT diff1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 1360
box 0 0 576 240
use JNWATR_PCH_4C1F2 diff1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 1600
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT diff1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 1360
box 0 0 576 240
use JNWATR_PCH_4C5F0 mirror1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 2000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP mirror1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 2400
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror3_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 0
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror3_MN4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 -240
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror4_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror4_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1088 0 1 800
box 0 0 576 240
use JNWATR_PCH_4C5F0 mirror1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP mirror1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2400
box 0 0 576 240
use JNWATR_PCH_12C5F0 mirror1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 3200
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP mirror1_MP3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 3600
box 0 0 832 240
use JNWATR_PCH_12CTAPBOT mirror1_MP3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 2960
box 0 0 832 240
use JNWATR_NCH_4C5F0 mirror4_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 400
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror4_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 800
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror3_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 0
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror3_MN3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1664 0 1 -240
box 0 0 576 240
use JNWATR_PCH_12C5F0 mirror1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 3200
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP mirror1_MP4_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 3600
box 0 0 832 240
use JNWATR_PCH_12CTAPBOT mirror1_MP4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 832 0 1 2960
box 0 0 832 240
use JNWTR_RPPO2 None_R1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 2496 0 1 0
box 0 0 724 1720
use JNWTR_RPPO2 None_R2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 0 0 1 0
box 0 0 724 1720
<< m1 >>
rect 1417 2013 1527 2067
<< m2 >>
rect 1417 2013 1527 2067
<< via1 >>
rect 1424 2020 1520 2060
<< m1 >>
rect 1417 13 1527 67
<< m2 >>
rect 1417 13 1527 67
<< via1 >>
rect 1424 20 1520 60
<< m1 >>
rect 1993 1613 2103 1667
<< m2 >>
rect 1993 1613 2103 1667
<< m3 >>
rect 1993 1613 2103 1667
<< via2 >>
rect 2000 1620 2096 1660
<< via1 >>
rect 2000 1620 2096 1660
<< m1 >>
rect 1161 173 1207 227
<< m2 >>
rect 1161 173 1207 227
<< via1 >>
rect 1168 180 1200 220
<< m1 >>
rect 1737 173 1783 227
<< m2 >>
rect 1737 173 1783 227
<< via1 >>
rect 1744 180 1776 220
<< m1 >>
rect 1993 13 2103 67
<< m2 >>
rect 1993 13 2103 67
<< via1 >>
rect 2000 20 2096 60
<< m1 >>
rect 1993 13 2103 67
<< m2 >>
rect 1993 13 2103 67
<< m3 >>
rect 1993 13 2103 67
<< via2 >>
rect 2000 20 2096 60
<< via1 >>
rect 2000 20 2096 60
<< m1 >>
rect 1801 1893 1911 1947
<< m2 >>
rect 1801 1893 1911 1947
<< via1 >>
rect 1808 1900 1904 1940
<< m1 >>
rect 1225 1893 1335 1947
<< m2 >>
rect 1225 1893 1335 1947
<< via1 >>
rect 1232 1900 1328 1940
<< m1 >>
rect 1417 3213 1527 3267
<< m2 >>
rect 1417 3213 1527 3267
<< via1 >>
rect 1424 3220 1520 3260
<< m1 >>
rect 1417 1613 1527 1667
<< m2 >>
rect 1417 1613 1527 1667
<< m3 >>
rect 1417 1613 1527 1667
<< via2 >>
rect 1424 1620 1520 1660
<< via1 >>
rect 1424 1620 1520 1660
<< m1 >>
rect 1161 573 1207 627
<< m2 >>
rect 1161 573 1207 627
<< via1 >>
rect 1168 580 1200 620
<< m1 >>
rect 1737 573 1783 627
<< m2 >>
rect 1737 573 1783 627
<< via1 >>
rect 1744 580 1776 620
<< m1 >>
rect 1161 2173 1207 2227
<< m2 >>
rect 1161 2173 1207 2227
<< via1 >>
rect 1168 2180 1200 2220
<< m1 >>
rect 1417 413 1527 467
<< m2 >>
rect 1417 413 1527 467
<< via1 >>
rect 1424 420 1520 460
<< m1 >>
rect 1737 2173 1783 2227
<< m2 >>
rect 1737 2173 1783 2227
<< via1 >>
rect 1744 2180 1776 2220
<< m1 >>
rect 1737 3373 1783 3427
<< m2 >>
rect 1737 3373 1783 3427
<< via1 >>
rect 1744 3380 1776 3420
<< m1 >>
rect 905 3373 951 3427
<< m2 >>
rect 905 3373 951 3427
<< via1 >>
rect 912 3380 944 3420
<< m1 >>
rect -250 3950 3470 4050
<< m1 >>
rect -250 -450 3470 -350
<< m1 >>
rect -250 -350 -150 3950
<< m1 >>
rect 3370 -350 3470 3950
<< m1 >>
rect -400 4100 3620 4200
<< m1 >>
rect -400 -600 3620 -500
<< m1 >>
rect -400 -500 -300 4100
<< m1 >>
rect 3520 -500 3620 4100
<< m2 >>
rect -213 2019 1466 2049
<< m3 >>
rect -213 19 -183 2049
<< m2 >>
rect -213 19 1466 49
<< m1 >>
rect 1417 2013 1527 2067
<< m2 >>
rect 1417 2013 1527 2067
<< via1 >>
rect 1424 2020 1520 2060
<< m1 >>
rect 1417 13 1527 67
<< m2 >>
rect 1417 13 1527 67
<< via1 >>
rect 1424 20 1520 60
<< m2 >>
rect -220 2012 -176 2056
<< m3 >>
rect -220 2012 -176 2056
<< via2 >>
rect -213 2019 -183 2049
<< m2 >>
rect -220 12 -176 56
<< m3 >>
rect -220 12 -176 56
<< via2 >>
rect -213 19 -183 49
<< m3 >>
rect 2030 822 2060 1637
<< m2 >>
rect 2030 822 2508 852
<< m3 >>
rect 2478 22 2508 852
<< m2 >>
rect 2030 22 2508 52
<< m3 >>
rect 2030 -410 2060 52
<< m2 >>
rect 2030 -410 2492 -380
<< m3 >>
rect 2462 -410 2492 212
<< m2 >>
rect 1181 182 2492 212
<< m1 >>
rect 1993 1613 2103 1667
<< m2 >>
rect 1993 1613 2103 1667
<< via1 >>
rect 2000 1620 2096 1660
<< m1 >>
rect 1161 173 1207 227
<< m2 >>
rect 1161 173 1207 227
<< via1 >>
rect 1168 180 1200 220
<< m1 >>
rect 1737 173 1783 227
<< m2 >>
rect 1737 173 1783 227
<< via1 >>
rect 1744 180 1776 220
<< m1 >>
rect 1993 13 2103 67
<< m2 >>
rect 1993 13 2103 67
<< via1 >>
rect 2000 20 2096 60
<< m1 >>
rect 1993 13 2103 67
<< m2 >>
rect 1993 13 2103 67
<< via1 >>
rect 2000 20 2096 60
<< m2 >>
rect 2023 815 2067 859
<< m3 >>
rect 2023 815 2067 859
<< via2 >>
rect 2030 822 2060 852
<< m2 >>
rect 2471 815 2515 859
<< m3 >>
rect 2471 815 2515 859
<< via2 >>
rect 2478 822 2508 852
<< m2 >>
rect 2471 15 2515 59
<< m3 >>
rect 2471 15 2515 59
<< via2 >>
rect 2478 22 2508 52
<< m2 >>
rect 2023 15 2067 59
<< m3 >>
rect 2023 15 2067 59
<< via2 >>
rect 2030 22 2060 52
<< m2 >>
rect 2023 -417 2067 -373
<< m3 >>
rect 2023 -417 2067 -373
<< via2 >>
rect 2030 -410 2060 -380
<< m2 >>
rect 2455 -417 2499 -373
<< m3 >>
rect 2455 -417 2499 -373
<< via2 >>
rect 2462 -410 2492 -380
<< m2 >>
rect 2455 175 2499 219
<< m3 >>
rect 2455 175 2499 219
<< via2 >>
rect 2462 182 2492 212
<< m2 >>
rect 813 1903 1852 1933
<< m3 >>
rect 813 1903 843 3245
<< m2 >>
rect 813 3215 1468 3245
<< m1 >>
rect 1801 1893 1911 1947
<< m2 >>
rect 1801 1893 1911 1947
<< via1 >>
rect 1808 1900 1904 1940
<< m1 >>
rect 1225 1893 1335 1947
<< m2 >>
rect 1225 1893 1335 1947
<< via1 >>
rect 1232 1900 1328 1940
<< m1 >>
rect 1417 3213 1527 3267
<< m2 >>
rect 1417 3213 1527 3267
<< via1 >>
rect 1424 3220 1520 3260
<< m2 >>
rect 806 1896 850 1940
<< m3 >>
rect 806 1896 850 1940
<< via2 >>
rect 813 1903 843 1933
<< m2 >>
rect 806 3208 850 3252
<< m3 >>
rect 806 3208 850 3252
<< via2 >>
rect 813 3215 843 3245
<< m3 >>
rect 1453 1189 1483 1636
<< m2 >>
rect 733 1189 1483 1219
<< m3 >>
rect 733 581 763 1219
<< m2 >>
rect 733 581 1756 611
<< m1 >>
rect 1417 1613 1527 1667
<< m2 >>
rect 1417 1613 1527 1667
<< via1 >>
rect 1424 1620 1520 1660
<< m1 >>
rect 1161 573 1207 627
<< m2 >>
rect 1161 573 1207 627
<< via1 >>
rect 1168 580 1200 620
<< m1 >>
rect 1737 573 1783 627
<< m2 >>
rect 1737 573 1783 627
<< via1 >>
rect 1744 580 1776 620
<< m2 >>
rect 1446 1182 1490 1226
<< m3 >>
rect 1446 1182 1490 1226
<< via2 >>
rect 1453 1189 1483 1219
<< m2 >>
rect 726 1182 770 1226
<< m3 >>
rect 726 1182 770 1226
<< via2 >>
rect 733 1189 763 1219
<< m2 >>
rect 726 574 770 618
<< m3 >>
rect 726 574 770 618
<< via2 >>
rect 733 581 763 611
<< m2 >>
rect 1180 2181 2315 2211
<< m3 >>
rect 2285 2181 2315 2643
<< m2 >>
rect 573 2613 2315 2643
<< m3 >>
rect 573 1621 603 2643
<< m2 >>
rect 573 1621 1035 1651
<< m3 >>
rect 1005 1093 1035 1651
<< m2 >>
rect 573 1093 1035 1123
<< m3 >>
rect 573 421 603 1123
<< m2 >>
rect 573 421 1468 451
<< m1 >>
rect 1161 2173 1207 2227
<< m2 >>
rect 1161 2173 1207 2227
<< via1 >>
rect 1168 2180 1200 2220
<< m1 >>
rect 1417 413 1527 467
<< m2 >>
rect 1417 413 1527 467
<< via1 >>
rect 1424 420 1520 460
<< m1 >>
rect 1737 2173 1783 2227
<< m2 >>
rect 1737 2173 1783 2227
<< via1 >>
rect 1744 2180 1776 2220
<< m2 >>
rect 2278 2174 2322 2218
<< m3 >>
rect 2278 2174 2322 2218
<< via2 >>
rect 2285 2181 2315 2211
<< m2 >>
rect 2278 2606 2322 2650
<< m3 >>
rect 2278 2606 2322 2650
<< via2 >>
rect 2285 2613 2315 2643
<< m2 >>
rect 566 2606 610 2650
<< m3 >>
rect 566 2606 610 2650
<< via2 >>
rect 573 2613 603 2643
<< m2 >>
rect 566 1614 610 1658
<< m3 >>
rect 566 1614 610 1658
<< via2 >>
rect 573 1621 603 1651
<< m2 >>
rect 998 1614 1042 1658
<< m3 >>
rect 998 1614 1042 1658
<< via2 >>
rect 1005 1621 1035 1651
<< m2 >>
rect 998 1086 1042 1130
<< m3 >>
rect 998 1086 1042 1130
<< via2 >>
rect 1005 1093 1035 1123
<< m2 >>
rect 566 1086 610 1130
<< m3 >>
rect 566 1086 610 1130
<< via2 >>
rect 573 1093 603 1123
<< m2 >>
rect 566 414 610 458
<< m3 >>
rect 566 414 610 458
<< via2 >>
rect 573 421 603 451
<< m2 >>
rect 922 3379 1754 3409
<< m1 >>
rect 1737 3373 1783 3427
<< m2 >>
rect 1737 3373 1783 3427
<< via1 >>
rect 1744 3380 1776 3420
<< m1 >>
rect 905 3373 951 3427
<< m2 >>
rect 905 3373 951 3427
<< via1 >>
rect 912 3380 944 3420
<< locali >>
rect 1040 2300 1328 2340
<< locali >>
rect 1040 300 1328 340
<< locali >>
rect 1040 700 1328 740
<< locali >>
rect 1616 2300 1904 2340
<< locali >>
rect 2000 2180 2160 2220
<< locali >>
rect 1616 3500 1904 3540
<< locali >>
rect 2256 3380 2416 3420
<< locali >>
rect 1616 700 1904 740
<< locali >>
rect 2000 580 2160 620
<< locali >>
rect 1616 300 1904 340
<< locali >>
rect 2000 180 2160 220
<< locali >>
rect 784 3500 1072 3540
<< locali >>
rect -250 1432 3470 1528
<< locali >>
rect -257 1425 -143 1535
<< m1 >>
rect -257 1425 -143 1535
<< viali >>
rect -250 1432 -150 1528
<< locali >>
rect 3363 1425 3477 1535
<< m1 >>
rect 3363 1425 3477 1535
<< viali >>
rect 3370 1432 3470 1528
<< locali >>
rect -250 2472 3470 2568
<< locali >>
rect -257 2465 -143 2575
<< m1 >>
rect -257 2465 -143 2575
<< viali >>
rect -250 2472 -150 2568
<< locali >>
rect 3363 2465 3477 2575
<< m1 >>
rect 3363 2465 3477 2575
<< viali >>
rect 3370 2472 3470 2568
<< locali >>
rect -400 -168 3620 -72
<< locali >>
rect -407 -175 -293 -65
<< m1 >>
rect -407 -175 -293 -65
<< viali >>
rect -400 -168 -300 -72
<< locali >>
rect 3513 -175 3627 -65
<< m1 >>
rect 3513 -175 3627 -65
<< viali >>
rect 3520 -168 3620 -72
<< locali >>
rect -400 872 3620 968
<< locali >>
rect -407 865 -293 975
<< m1 >>
rect -407 865 -293 975
<< viali >>
rect -400 872 -300 968
<< locali >>
rect 3513 865 3627 975
<< m1 >>
rect 3513 865 3627 975
<< viali >>
rect 3520 872 3620 968
<< locali >>
rect -250 3672 3470 3768
<< locali >>
rect -257 3665 -143 3775
<< m1 >>
rect -257 3665 -143 3775
<< viali >>
rect -250 3672 -150 3768
<< locali >>
rect 3363 3665 3477 3775
<< m1 >>
rect 3363 3665 3477 3775
<< viali >>
rect 3370 3672 3470 3768
<< locali >>
rect -250 3032 3470 3128
<< locali >>
rect -257 3025 -143 3135
<< m1 >>
rect -257 3025 -143 3135
<< viali >>
rect -250 3032 -150 3128
<< locali >>
rect 3363 3025 3477 3135
<< m1 >>
rect 3363 3025 3477 3135
<< viali >>
rect 3370 3032 3470 3128
<< locali >>
rect -250 3672 3470 3768
<< locali >>
rect -257 3665 -143 3775
<< m1 >>
rect -257 3665 -143 3775
<< viali >>
rect -250 3672 -150 3768
<< locali >>
rect 3363 3665 3477 3775
<< m1 >>
rect 3363 3665 3477 3775
<< viali >>
rect 3370 3672 3470 3768
<< labels >>
flabel m1 s -250 3950 3470 4050 0 FreeSans 400 0 0 0 VDD
port 1 nsew signal bidirectional
flabel m1 s -400 4100 3620 4200 0 FreeSans 400 0 0 0 VSS
port 2 nsew signal bidirectional
flabel m1 s 1168 1780 1200 1820 0 FreeSans 400 0 0 0 V_n
port 3 nsew signal bidirectional
flabel m1 s 1744 1780 1776 1820 0 FreeSans 400 0 0 0 V_p
port 4 nsew signal bidirectional
flabel m2 s -213 2019 1466 2049 0 FreeSans 400 0 0 0 I_out
port 5 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1745323676
<< checkpaint >>
rect 0 0 1000 1000
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 8960
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 8720
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8960
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8720
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 9360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9360
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 10160
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 10160
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 9760
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 9760
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 10560
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 10960
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 10560
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 10960
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 7760
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 8160
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 7520
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 7760
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 8160
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 7520
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 500
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 5340
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 300 0 1 2920
box 0 0 2236 1720
<< locali >>
rect 100 11310 2736 11360
<< locali >>
rect 100 100 2736 150
<< m1 >>
rect 100 150 150 11310
<< m1 >>
rect 2686 150 2736 11310
<< locali >>
rect 93 11303 157 11367
<< m1 >>
rect 93 11303 157 11367
<< viali >>
rect 100 11310 150 11360
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2679 11303 2743 11367
<< m1 >>
rect 2679 11303 2743 11367
<< viali >>
rect 2686 11310 2736 11360
<< locali >>
rect 2679 93 2743 157
<< m1 >>
rect 2679 93 2743 157
<< viali >>
rect 2686 100 2736 150
<< locali >>
rect 0 11410 2836 11460
<< locali >>
rect 0 0 2836 50
<< m1 >>
rect 0 50 50 11410
<< m1 >>
rect 2786 50 2836 11410
<< locali >>
rect -7 11403 57 11467
<< m1 >>
rect -7 11403 57 11467
<< viali >>
rect 0 11410 50 11460
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2779 11403 2843 11467
<< m1 >>
rect 2779 11403 2843 11467
<< viali >>
rect 2786 11410 2836 11460
<< locali >>
rect 2779 -7 2843 57
<< m1 >>
rect 2779 -7 2843 57
<< viali >>
rect 2786 0 2836 50
<< locali >>
rect 252 10860 540 10900
<< locali >>
rect 828 10860 1116 10900
<< locali >>
rect 1212 10740 1372 10780
<< locali >>
rect 252 8060 540 8100
<< locali >>
rect 636 7940 796 7980
<< locali >>
rect 828 8060 1116 8100
<< locali >>
rect 100 8792 2736 8888
<< locali >>
rect 93 8785 157 8895
<< m1 >>
rect 93 8785 157 8895
<< viali >>
rect 100 8792 150 8888
<< locali >>
rect 2679 8785 2743 8895
<< m1 >>
rect 2679 8785 2743 8895
<< viali >>
rect 2686 8792 2736 8888
<< locali >>
rect 100 11032 2736 11128
<< locali >>
rect 93 11025 157 11135
<< m1 >>
rect 93 11025 157 11135
<< viali >>
rect 100 11032 150 11128
<< locali >>
rect 2679 11025 2743 11135
<< m1 >>
rect 2679 11025 2743 11135
<< viali >>
rect 2686 11032 2736 11128
<< locali >>
rect 0 8232 2836 8328
<< locali >>
rect -7 8225 57 8335
<< m1 >>
rect -7 8225 57 8335
<< viali >>
rect 0 8232 50 8328
<< locali >>
rect 2779 8225 2843 8335
<< m1 >>
rect 2779 8225 2843 8335
<< viali >>
rect 2786 8232 2836 8328
<< locali >>
rect 0 7592 2836 7688
<< locali >>
rect -7 7585 57 7695
<< m1 >>
rect -7 7585 57 7695
<< viali >>
rect 0 7592 50 7688
<< locali >>
rect 2779 7585 2843 7695
<< m1 >>
rect 2779 7585 2843 7695
<< viali >>
rect 2786 7592 2836 7688
<< labels >>
flabel locali s 100 11310 2736 11360 0 FreeSans 400 0 0 0 VDD
port 78 nsew signal bidirectional
flabel locali s 0 11410 2836 11460 0 FreeSans 400 0 0 0 VSS
port 79 nsew signal bidirectional
<< properties >>
<< end >>
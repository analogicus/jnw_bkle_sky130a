magic
tech sky130A
magscale 1 1
timestamp 1740580848
<< checkpaint >>
rect 0 0 0 0
use COMP COMP 
transform 1 0 0 0 1 0
box 1674 50 2826 3850
<< labels >>
<< properties >>
<< end >>
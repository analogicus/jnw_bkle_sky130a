magic
tech sky130A
magscale 1 1
timestamp 1737386094
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 MN1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 1500
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN2 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 1500
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP5 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 100
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP6 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 100
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 900
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP2 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 900
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN3 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 2300
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN4 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 2300
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN5 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 1900
box 0 0 576 400
use JNWATR_NCH_4C5F0 MN6 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 1900
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP3 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 924 0 1 500
box 0 0 576 400
use JNWATR_PCH_4C5F0 MP4 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_COMP_LIBS/JNW_ATR_SKY130A
transform 1 0 1500 0 1 500
box 0 0 576 400
<< m1 >>
rect 1061 1793 1171 1847
<< m2 >>
rect 1061 1793 1171 1847
<< m3 >>
rect 1061 1793 1171 1847
<< via2 >>
rect 1068 1800 1164 1840
<< via1 >>
rect 1068 1800 1164 1840
<< locali >>
rect 869 1673 979 1727
<< m1 >>
rect 869 1673 979 1727
<< m2 >>
rect 869 1673 979 1727
<< via1 >>
rect 876 1680 972 1720
<< viali >>
rect 876 1680 972 1720
<< m1 >>
rect 1637 1793 1747 1847
<< m2 >>
rect 1637 1793 1747 1847
<< m3 >>
rect 1637 1793 1747 1847
<< via2 >>
rect 1644 1800 1740 1840
<< via1 >>
rect 1644 1800 1740 1840
<< locali >>
rect 1445 1673 1555 1727
<< m1 >>
rect 1445 1673 1555 1727
<< m2 >>
rect 1445 1673 1555 1727
<< via1 >>
rect 1452 1680 1548 1720
<< viali >>
rect 1452 1680 1548 1720
<< m1 >>
rect 1061 393 1171 447
<< m2 >>
rect 1061 393 1171 447
<< m3 >>
rect 1061 393 1171 447
<< via2 >>
rect 1068 400 1164 440
<< via1 >>
rect 1068 400 1164 440
<< locali >>
rect 869 273 979 327
<< m1 >>
rect 869 273 979 327
<< m2 >>
rect 869 273 979 327
<< via1 >>
rect 876 280 972 320
<< viali >>
rect 876 280 972 320
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< m3 >>
rect 1637 393 1747 447
<< via2 >>
rect 1644 400 1740 440
<< via1 >>
rect 1644 400 1740 440
<< locali >>
rect 1445 273 1555 327
<< m1 >>
rect 1445 273 1555 327
<< m2 >>
rect 1445 273 1555 327
<< via1 >>
rect 1452 280 1548 320
<< viali >>
rect 1452 280 1548 320
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< locali >>
rect 869 1073 979 1127
<< m1 >>
rect 869 1073 979 1127
<< m2 >>
rect 869 1073 979 1127
<< via1 >>
rect 876 1080 972 1120
<< viali >>
rect 876 1080 972 1120
<< m1 >>
rect 1573 1073 1619 1127
<< m2 >>
rect 1573 1073 1619 1127
<< via1 >>
rect 1580 1080 1612 1120
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< m3 >>
rect 1829 913 1939 967
<< via2 >>
rect 1836 920 1932 960
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< m1 >>
rect 1061 2593 1171 2647
<< m2 >>
rect 1061 2593 1171 2647
<< m3 >>
rect 1061 2593 1171 2647
<< via2 >>
rect 1068 2600 1164 2640
<< via1 >>
rect 1068 2600 1164 2640
<< locali >>
rect 869 2473 979 2527
<< m1 >>
rect 869 2473 979 2527
<< m2 >>
rect 869 2473 979 2527
<< via1 >>
rect 876 2480 972 2520
<< viali >>
rect 876 2480 972 2520
<< m1 >>
rect 1573 2473 1619 2527
<< m2 >>
rect 1573 2473 1619 2527
<< via1 >>
rect 1580 2480 1612 2520
<< m1 >>
rect 1829 2313 1939 2367
<< m2 >>
rect 1829 2313 1939 2367
<< m3 >>
rect 1829 2313 1939 2367
<< via2 >>
rect 1836 2320 1932 2360
<< via1 >>
rect 1836 2320 1932 2360
<< m1 >>
rect 1637 2593 1747 2647
<< m2 >>
rect 1637 2593 1747 2647
<< m3 >>
rect 1637 2593 1747 2647
<< via2 >>
rect 1644 2600 1740 2640
<< via1 >>
rect 1644 2600 1740 2640
<< locali >>
rect 1445 2473 1555 2527
<< m1 >>
rect 1445 2473 1555 2527
<< m2 >>
rect 1445 2473 1555 2527
<< via1 >>
rect 1452 2480 1548 2520
<< viali >>
rect 1452 2480 1548 2520
<< m1 >>
rect 997 2073 1043 2127
<< m2 >>
rect 997 2073 1043 2127
<< via1 >>
rect 1004 2080 1036 2120
<< m1 >>
rect 1253 1913 1363 1967
<< m2 >>
rect 1253 1913 1363 1967
<< m3 >>
rect 1253 1913 1363 1967
<< via2 >>
rect 1260 1920 1356 1960
<< via1 >>
rect 1260 1920 1356 1960
<< m1 >>
rect 1061 2193 1171 2247
<< m2 >>
rect 1061 2193 1171 2247
<< m3 >>
rect 1061 2193 1171 2247
<< via2 >>
rect 1068 2200 1164 2240
<< via1 >>
rect 1068 2200 1164 2240
<< locali >>
rect 869 2073 979 2127
<< m1 >>
rect 869 2073 979 2127
<< m2 >>
rect 869 2073 979 2127
<< via1 >>
rect 876 2080 972 2120
<< viali >>
rect 876 2080 972 2120
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< m3 >>
rect 1637 2193 1747 2247
<< via2 >>
rect 1644 2200 1740 2240
<< via1 >>
rect 1644 2200 1740 2240
<< locali >>
rect 1445 2073 1555 2127
<< m1 >>
rect 1445 2073 1555 2127
<< m2 >>
rect 1445 2073 1555 2127
<< via1 >>
rect 1452 2080 1548 2120
<< viali >>
rect 1452 2080 1548 2120
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< m3 >>
rect 1061 793 1171 847
<< via2 >>
rect 1068 800 1164 840
<< via1 >>
rect 1068 800 1164 840
<< locali >>
rect 869 673 979 727
<< m1 >>
rect 869 673 979 727
<< m2 >>
rect 869 673 979 727
<< via1 >>
rect 876 680 972 720
<< viali >>
rect 876 680 972 720
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1829 1513 1939 1567
<< m2 >>
rect 1829 1513 1939 1567
<< via1 >>
rect 1836 1520 1932 1560
<< m1 >>
rect 1829 113 1939 167
<< m2 >>
rect 1829 113 1939 167
<< via1 >>
rect 1836 120 1932 160
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1829 1913 1939 1967
<< m2 >>
rect 1829 1913 1939 1967
<< via1 >>
rect 1836 1920 1932 1960
<< m1 >>
rect 1829 1913 1939 1967
<< m2 >>
rect 1829 1913 1939 1967
<< via1 >>
rect 1836 1920 1932 1960
<< m1 >>
rect 1829 513 1939 567
<< m2 >>
rect 1829 513 1939 567
<< via1 >>
rect 1836 520 1932 560
<< m1 >>
rect 1573 273 1619 327
<< m2 >>
rect 1573 273 1619 327
<< via1 >>
rect 1580 280 1612 320
<< m1 >>
rect 997 673 1043 727
<< m2 >>
rect 997 673 1043 727
<< via1 >>
rect 1004 680 1036 720
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1573 273 1619 327
<< m2 >>
rect 1573 273 1619 327
<< m3 >>
rect 1573 273 1619 327
<< via2 >>
rect 1580 280 1612 320
<< via1 >>
rect 1580 280 1612 320
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1829 513 1939 567
<< m2 >>
rect 1829 513 1939 567
<< m3 >>
rect 1829 513 1939 567
<< via2 >>
rect 1836 520 1932 560
<< via1 >>
rect 1836 520 1932 560
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 393 1747 447
<< m2 >>
rect 1637 393 1747 447
<< via1 >>
rect 1644 400 1740 440
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 997 1073 1043 1127
<< m2 >>
rect 997 1073 1043 1127
<< via1 >>
rect 1004 1080 1036 1120
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< m3 >>
rect 1061 1193 1171 1247
<< via2 >>
rect 1068 1200 1164 1240
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< m3 >>
rect 1637 1193 1747 1247
<< via2 >>
rect 1644 1200 1740 1240
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1637 1193 1747 1247
<< m2 >>
rect 1637 1193 1747 1247
<< via1 >>
rect 1644 1200 1740 1240
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1253 1913 1363 1967
<< m2 >>
rect 1253 1913 1363 1967
<< via1 >>
rect 1260 1920 1356 1960
<< m1 >>
rect 1253 1913 1363 1967
<< m2 >>
rect 1253 1913 1363 1967
<< via1 >>
rect 1260 1920 1356 1960
<< m1 >>
rect 1253 1513 1363 1567
<< m2 >>
rect 1253 1513 1363 1567
<< via1 >>
rect 1260 1520 1356 1560
<< m1 >>
rect 1253 913 1363 967
<< m2 >>
rect 1253 913 1363 967
<< via1 >>
rect 1260 920 1356 960
<< m1 >>
rect 1253 1913 1363 1967
<< m2 >>
rect 1253 1913 1363 1967
<< via1 >>
rect 1260 1920 1356 1960
<< m1 >>
rect 1573 2073 1619 2127
<< m2 >>
rect 1573 2073 1619 2127
<< m3 >>
rect 1573 2073 1619 2127
<< via2 >>
rect 1580 2080 1612 2120
<< via1 >>
rect 1580 2080 1612 2120
<< locali >>
rect 1445 2073 1555 2127
<< m1 >>
rect 1445 2073 1555 2127
<< m2 >>
rect 1445 2073 1555 2127
<< via1 >>
rect 1452 2080 1548 2120
<< viali >>
rect 1452 2080 1548 2120
<< locali >>
rect 1445 2073 1555 2127
<< m1 >>
rect 1445 2073 1555 2127
<< m2 >>
rect 1445 2073 1555 2127
<< m3 >>
rect 1445 2073 1555 2127
<< via2 >>
rect 1452 2080 1548 2120
<< via1 >>
rect 1452 2080 1548 2120
<< viali >>
rect 1452 2080 1548 2120
<< m1 >>
rect 997 1073 1043 1127
<< m2 >>
rect 997 1073 1043 1127
<< m3 >>
rect 997 1073 1043 1127
<< via2 >>
rect 1004 1080 1036 1120
<< via1 >>
rect 1004 1080 1036 1120
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< m3 >>
rect 1253 513 1363 567
<< via2 >>
rect 1260 520 1356 560
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 1061 793 1171 847
<< m2 >>
rect 1061 793 1171 847
<< via1 >>
rect 1068 800 1164 840
<< m1 >>
rect 997 1073 1043 1127
<< m2 >>
rect 997 1073 1043 1127
<< m3 >>
rect 997 1073 1043 1127
<< via2 >>
rect 1004 1080 1036 1120
<< via1 >>
rect 1004 1080 1036 1120
<< m1 >>
rect 1573 673 1619 727
<< m2 >>
rect 1573 673 1619 727
<< m3 >>
rect 1573 673 1619 727
<< via2 >>
rect 1580 680 1612 720
<< via1 >>
rect 1580 680 1612 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 1061 1193 1171 1247
<< m2 >>
rect 1061 1193 1171 1247
<< via1 >>
rect 1068 1200 1164 1240
<< locali >>
rect 1445 1073 1555 1127
<< m1 >>
rect 1445 1073 1555 1127
<< m2 >>
rect 1445 1073 1555 1127
<< via1 >>
rect 1452 1080 1548 1120
<< viali >>
rect 1452 1080 1548 1120
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1253 513 1363 567
<< m2 >>
rect 1253 513 1363 567
<< via1 >>
rect 1260 520 1356 560
<< m1 >>
rect 1573 673 1619 727
<< m2 >>
rect 1573 673 1619 727
<< m3 >>
rect 1573 673 1619 727
<< via2 >>
rect 1580 680 1612 720
<< via1 >>
rect 1580 680 1612 720
<< locali >>
rect 1445 673 1555 727
<< m1 >>
rect 1445 673 1555 727
<< m2 >>
rect 1445 673 1555 727
<< m3 >>
rect 1445 673 1555 727
<< via2 >>
rect 1452 680 1548 720
<< via1 >>
rect 1452 680 1548 720
<< viali >>
rect 1452 680 1548 720
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< m3 >>
rect 1829 913 1939 967
<< via2 >>
rect 1836 920 1932 960
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1829 913 1939 967
<< m2 >>
rect 1829 913 1939 967
<< via1 >>
rect 1836 920 1932 960
<< m1 >>
rect 1573 673 1619 727
<< m2 >>
rect 1573 673 1619 727
<< via1 >>
rect 1580 680 1612 720
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< m3 >>
rect 1637 793 1747 847
<< via2 >>
rect 1644 800 1740 840
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 1637 793 1747 847
<< m2 >>
rect 1637 793 1747 847
<< via1 >>
rect 1644 800 1740 840
<< m1 >>
rect 997 2473 1043 2527
<< m2 >>
rect 997 2473 1043 2527
<< via1 >>
rect 1004 2480 1036 2520
<< m1 >>
rect 1829 2313 1939 2367
<< m2 >>
rect 1829 2313 1939 2367
<< via1 >>
rect 1836 2320 1932 2360
<< m1 >>
rect 1829 2313 1939 2367
<< m2 >>
rect 1829 2313 1939 2367
<< m3 >>
rect 1829 2313 1939 2367
<< via2 >>
rect 1836 2320 1932 2360
<< via1 >>
rect 1836 2320 1932 2360
<< m1 >>
rect 1061 2593 1171 2647
<< m2 >>
rect 1061 2593 1171 2647
<< m3 >>
rect 1061 2593 1171 2647
<< via2 >>
rect 1068 2600 1164 2640
<< via1 >>
rect 1068 2600 1164 2640
<< m1 >>
rect 1637 2593 1747 2647
<< m2 >>
rect 1637 2593 1747 2647
<< m3 >>
rect 1637 2593 1747 2647
<< via2 >>
rect 1644 2600 1740 2640
<< via1 >>
rect 1644 2600 1740 2640
<< m1 >>
rect 1061 2593 1171 2647
<< m2 >>
rect 1061 2593 1171 2647
<< via1 >>
rect 1068 2600 1164 2640
<< m1 >>
rect 1061 2193 1171 2247
<< m2 >>
rect 1061 2193 1171 2247
<< via1 >>
rect 1068 2200 1164 2240
<< m1 >>
rect 1061 2593 1171 2647
<< m2 >>
rect 1061 2593 1171 2647
<< m3 >>
rect 1061 2593 1171 2647
<< via2 >>
rect 1068 2600 1164 2640
<< via1 >>
rect 1068 2600 1164 2640
<< m1 >>
rect 1061 2593 1171 2647
<< m2 >>
rect 1061 2593 1171 2647
<< via1 >>
rect 1068 2600 1164 2640
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< via1 >>
rect 1644 2200 1740 2240
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< m3 >>
rect 1637 2193 1747 2247
<< via2 >>
rect 1644 2200 1740 2240
<< via1 >>
rect 1644 2200 1740 2240
<< m1 >>
rect 1573 2473 1619 2527
<< m2 >>
rect 1573 2473 1619 2527
<< m3 >>
rect 1573 2473 1619 2527
<< via2 >>
rect 1580 2480 1612 2520
<< via1 >>
rect 1580 2480 1612 2520
<< m1 >>
rect 1637 2593 1747 2647
<< m2 >>
rect 1637 2593 1747 2647
<< via1 >>
rect 1644 2600 1740 2640
<< locali >>
rect 1445 2473 1555 2527
<< m1 >>
rect 1445 2473 1555 2527
<< m2 >>
rect 1445 2473 1555 2527
<< m3 >>
rect 1445 2473 1555 2527
<< via2 >>
rect 1452 2480 1548 2520
<< via1 >>
rect 1452 2480 1548 2520
<< viali >>
rect 1452 2480 1548 2520
<< m1 >>
rect 1061 2193 1171 2247
<< m2 >>
rect 1061 2193 1171 2247
<< m3 >>
rect 1061 2193 1171 2247
<< via2 >>
rect 1068 2200 1164 2240
<< via1 >>
rect 1068 2200 1164 2240
<< m1 >>
rect 1637 2593 1747 2647
<< m2 >>
rect 1637 2593 1747 2647
<< via1 >>
rect 1644 2600 1740 2640
<< m1 >>
rect 1637 2593 1747 2647
<< m2 >>
rect 1637 2593 1747 2647
<< via1 >>
rect 1644 2600 1740 2640
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< via1 >>
rect 1644 2200 1740 2240
<< m1 >>
rect 1253 1913 1363 1967
<< m2 >>
rect 1253 1913 1363 1967
<< m3 >>
rect 1253 1913 1363 1967
<< via2 >>
rect 1260 1920 1356 1960
<< via1 >>
rect 1260 1920 1356 1960
<< m1 >>
rect 1573 2073 1619 2127
<< m2 >>
rect 1573 2073 1619 2127
<< via1 >>
rect 1580 2080 1612 2120
<< m1 >>
rect 1061 2193 1171 2247
<< m2 >>
rect 1061 2193 1171 2247
<< via1 >>
rect 1068 2200 1164 2240
<< m1 >>
rect 1061 2193 1171 2247
<< m2 >>
rect 1061 2193 1171 2247
<< m3 >>
rect 1061 2193 1171 2247
<< via2 >>
rect 1068 2200 1164 2240
<< via1 >>
rect 1068 2200 1164 2240
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< m3 >>
rect 1637 2193 1747 2247
<< via2 >>
rect 1644 2200 1740 2240
<< via1 >>
rect 1644 2200 1740 2240
<< m1 >>
rect 1637 2193 1747 2247
<< m2 >>
rect 1637 2193 1747 2247
<< via1 >>
rect 1644 2200 1740 2240
<< m1 >>
rect 997 673 1043 727
<< m2 >>
rect 997 673 1043 727
<< m3 >>
rect 997 673 1043 727
<< via2 >>
rect 1004 680 1036 720
<< via1 >>
rect 1004 680 1036 720
<< m1 >>
rect 1829 513 1939 567
<< m2 >>
rect 1829 513 1939 567
<< m3 >>
rect 1829 513 1939 567
<< via2 >>
rect 1836 520 1932 560
<< via1 >>
rect 1836 520 1932 560
<< m3 >>
rect 909 1805 1116 1835
<< m2 >>
rect 909 1700 939 1835
<< m2 >>
rect 902 1798 946 1842
<< m3 >>
rect 902 1798 946 1842
<< via2 >>
rect 909 1805 939 1835
<< m3 >>
rect 1500 1805 1692 1835
<< m2 >>
rect 1485 1700 1515 1820
<< m2 >>
rect 1493 1798 1522 1827
<< m3 >>
rect 1493 1798 1522 1827
<< via2 >>
rect 1500 1805 1515 1820
<< m3 >>
rect 924 405 1116 435
<< m2 >>
rect 909 300 939 420
<< m2 >>
rect 917 398 946 427
<< m3 >>
rect 917 398 946 427
<< via2 >>
rect 924 405 939 420
<< m3 >>
rect 1500 405 1692 435
<< m2 >>
rect 1485 300 1515 420
<< m2 >>
rect 1493 398 1522 427
<< m3 >>
rect 1493 398 1522 427
<< via2 >>
rect 1500 405 1515 420
<< m3 >>
rect 924 1205 1116 1235
<< m2 >>
rect 909 1100 939 1220
<< m2 >>
rect 917 1198 946 1227
<< m3 >>
rect 917 1198 946 1227
<< via2 >>
rect 924 1205 939 1220
<< m3 >>
rect 1596 925 1884 955
<< m2 >>
rect 1581 940 1611 1100
<< m2 >>
rect 1589 933 1618 962
<< m3 >>
rect 1589 933 1618 962
<< via2 >>
rect 1596 940 1611 955
<< m3 >>
rect 1500 1205 1692 1235
<< m2 >>
rect 1485 1100 1515 1220
<< m2 >>
rect 1493 1198 1522 1227
<< m3 >>
rect 1493 1198 1522 1227
<< via2 >>
rect 1500 1205 1515 1220
<< m3 >>
rect 924 2605 1116 2635
<< m2 >>
rect 909 2500 939 2620
<< m2 >>
rect 917 2598 946 2627
<< m3 >>
rect 917 2598 946 2627
<< via2 >>
rect 924 2605 939 2620
<< m3 >>
rect 1596 2325 1884 2355
<< m2 >>
rect 1581 2340 1611 2500
<< m2 >>
rect 1589 2333 1618 2362
<< m3 >>
rect 1589 2333 1618 2362
<< via2 >>
rect 1596 2340 1611 2355
<< m3 >>
rect 1500 2605 1692 2635
<< m2 >>
rect 1485 2500 1515 2620
<< m2 >>
rect 1493 2598 1522 2627
<< m3 >>
rect 1493 2598 1522 2627
<< via2 >>
rect 1500 2605 1515 2620
<< m3 >>
rect 1005 1925 1308 1955
<< m2 >>
rect 1005 1925 1035 2100
<< m2 >>
rect 998 1918 1042 1962
<< m3 >>
rect 998 1918 1042 1962
<< via2 >>
rect 1005 1925 1035 1955
<< m3 >>
rect 924 2205 1116 2235
<< m2 >>
rect 909 2100 939 2220
<< m2 >>
rect 917 2198 946 2227
<< m3 >>
rect 917 2198 946 2227
<< via2 >>
rect 924 2205 939 2220
<< m3 >>
rect 1485 2205 1692 2235
<< m2 >>
rect 1485 2100 1515 2235
<< m2 >>
rect 1478 2198 1522 2242
<< m3 >>
rect 1478 2198 1522 2242
<< via2 >>
rect 1485 2205 1515 2235
<< m3 >>
rect 924 805 1116 835
<< m2 >>
rect 909 700 939 820
<< m2 >>
rect 917 798 946 827
<< m3 >>
rect 917 798 946 827
<< via2 >>
rect 924 805 939 820
<< m3 >>
rect 1500 805 1692 835
<< m2 >>
rect 1485 700 1515 820
<< m2 >>
rect 1493 798 1522 827
<< m3 >>
rect 1493 798 1522 827
<< via2 >>
rect 1500 805 1515 820
<< m2 >>
rect 1677 420 1707 477
<< m3 >>
rect 1180 462 1692 492
<< m2 >>
rect 1165 477 1195 877
<< m3 >>
rect 1116 862 1180 892
<< m2 >>
rect 1101 877 1131 1220
<< m2 >>
rect 1670 455 1699 484
<< m3 >>
rect 1670 455 1699 484
<< via2 >>
rect 1677 462 1692 477
<< m2 >>
rect 1173 470 1202 499
<< m3 >>
rect 1173 470 1202 499
<< via2 >>
rect 1180 477 1195 492
<< m2 >>
rect 1158 855 1187 884
<< m3 >>
rect 1158 855 1187 884
<< via2 >>
rect 1165 862 1180 877
<< m2 >>
rect 1109 870 1138 899
<< m3 >>
rect 1109 870 1138 899
<< via2 >>
rect 1116 877 1131 892
<< m2 >>
rect 1677 420 1707 727
<< m2 >>
rect 1677 727 1707 727
<< m2 >>
rect 1677 727 1707 1220
<< m2 >>
rect 1677 1220 1707 1220
<< m2 >>
rect 1869 140 1899 388
<< m2 >>
rect 1869 388 1899 388
<< m2 >>
rect 1869 388 1899 1940
<< m2 >>
rect 1869 1940 1899 1940
<< m2 >>
rect 1581 300 1611 357
<< m3 >>
rect 1020 342 1596 372
<< m2 >>
rect 1005 357 1035 700
<< m2 >>
rect 1574 335 1603 364
<< m3 >>
rect 1574 335 1603 364
<< via2 >>
rect 1581 342 1596 357
<< m2 >>
rect 1013 350 1042 379
<< m3 >>
rect 1013 350 1042 379
<< via2 >>
rect 1020 357 1035 372
<< m2 >>
rect 1677 420 1707 464
<< m3 >>
rect 1628 449 1692 479
<< m2 >>
rect 1613 464 1643 597
<< m3 >>
rect 1372 582 1628 612
<< m2 >>
rect 1357 597 1387 642
<< m3 >>
rect 1116 627 1372 657
<< m2 >>
rect 1101 642 1131 820
<< m2 >>
rect 1670 442 1699 471
<< m3 >>
rect 1670 442 1699 471
<< via2 >>
rect 1677 449 1692 464
<< m2 >>
rect 1621 457 1650 486
<< m3 >>
rect 1621 457 1650 486
<< via2 >>
rect 1628 464 1643 479
<< m2 >>
rect 1606 575 1635 604
<< m3 >>
rect 1606 575 1635 604
<< via2 >>
rect 1613 582 1628 597
<< m2 >>
rect 1365 590 1394 619
<< m3 >>
rect 1365 590 1394 619
<< via2 >>
rect 1372 597 1387 612
<< m2 >>
rect 1350 620 1379 649
<< m3 >>
rect 1350 620 1379 649
<< via2 >>
rect 1357 627 1372 642
<< m2 >>
rect 1109 635 1138 664
<< m3 >>
rect 1109 635 1138 664
<< via2 >>
rect 1116 642 1131 657
<< m3 >>
rect 1596 285 1668 315
<< m2 >>
rect 1653 300 1683 360
<< m3 >>
rect 1668 345 1740 375
<< m2 >>
rect 1725 360 1755 540
<< m3 >>
rect 1740 525 1884 555
<< m2 >>
rect 1646 293 1675 322
<< m3 >>
rect 1646 293 1675 322
<< via2 >>
rect 1653 300 1668 315
<< m2 >>
rect 1661 338 1690 367
<< m3 >>
rect 1661 338 1690 367
<< via2 >>
rect 1668 345 1683 360
<< m2 >>
rect 1718 353 1747 382
<< m3 >>
rect 1718 353 1747 382
<< via2 >>
rect 1725 360 1740 375
<< m2 >>
rect 1733 518 1762 547
<< m3 >>
rect 1733 518 1762 547
<< via2 >>
rect 1740 525 1755 540
<< m2 >>
rect 1677 420 1707 420
<< m2 >>
rect 1677 420 1707 591
<< m2 >>
rect 1677 591 1707 591
<< m2 >>
rect 1677 591 1707 820
<< m2 >>
rect 1677 820 1707 820
<< m2 >>
rect 1005 1020 1035 1100
<< m3 >>
rect 1020 1005 1884 1035
<< m2 >>
rect 1869 940 1899 1020
<< m2 >>
rect 1013 1013 1042 1042
<< m3 >>
rect 1013 1013 1042 1042
<< via2 >>
rect 1020 1020 1035 1035
<< m2 >>
rect 1862 998 1891 1027
<< m3 >>
rect 1862 998 1891 1027
<< via2 >>
rect 1869 1005 1884 1020
<< m3 >>
rect 1116 1205 1372 1235
<< m2 >>
rect 1357 1220 1387 1220
<< m3 >>
rect 1372 1205 1692 1235
<< m2 >>
rect 1677 1220 1707 1220
<< m2 >>
rect 1293 940 1323 1440
<< m2 >>
rect 1293 1440 1323 1440
<< m2 >>
rect 1293 1440 1323 1940
<< m2 >>
rect 1293 1940 1323 1940
<< m2 >>
rect 1293 940 1323 1004
<< m3 >>
rect 1308 989 1365 1019
<< m2 >>
rect 1350 1004 1380 2035
<< m3 >>
rect 1365 2020 1538 2050
<< m2 >>
rect 1523 2035 1553 2100
<< m3 >>
rect 1538 2085 1596 2115
<< m2 >>
rect 1301 982 1330 1011
<< m3 >>
rect 1301 982 1330 1011
<< via2 >>
rect 1308 989 1323 1004
<< m2 >>
rect 1343 997 1372 1026
<< m3 >>
rect 1343 997 1372 1026
<< via2 >>
rect 1350 1004 1365 1019
<< m2 >>
rect 1358 2013 1387 2042
<< m3 >>
rect 1358 2013 1387 2042
<< via2 >>
rect 1365 2020 1380 2035
<< m2 >>
rect 1516 2028 1545 2057
<< m3 >>
rect 1516 2028 1545 2057
<< via2 >>
rect 1523 2035 1538 2050
<< m2 >>
rect 1531 2078 1560 2107
<< m3 >>
rect 1531 2078 1560 2107
<< via2 >>
rect 1538 2085 1553 2100
<< m3 >>
rect 1020 1085 1077 1115
<< m2 >>
rect 1062 540 1092 1100
<< m3 >>
rect 1077 525 1308 555
<< m2 >>
rect 1055 1078 1084 1107
<< m3 >>
rect 1055 1078 1084 1107
<< via2 >>
rect 1062 1085 1077 1100
<< m2 >>
rect 1070 533 1099 562
<< m3 >>
rect 1070 533 1099 562
<< via2 >>
rect 1077 540 1092 555
<< m2 >>
rect 1101 934 1131 1220
<< m2 >>
rect 1101 934 1131 934
<< m2 >>
rect 1101 820 1131 934
<< m2 >>
rect 1101 820 1131 820
<< m3 >>
rect 1020 1085 1404 1115
<< m2 >>
rect 1389 757 1419 1100
<< m3 >>
rect 1404 742 1532 772
<< m2 >>
rect 1517 700 1547 757
<< m3 >>
rect 1532 685 1596 715
<< m2 >>
rect 1382 1078 1411 1107
<< m3 >>
rect 1382 1078 1411 1107
<< via2 >>
rect 1389 1085 1404 1100
<< m2 >>
rect 1397 750 1426 779
<< m3 >>
rect 1397 750 1426 779
<< via2 >>
rect 1404 757 1419 772
<< m2 >>
rect 1510 735 1539 764
<< m3 >>
rect 1510 735 1539 764
<< via2 >>
rect 1517 742 1532 757
<< m2 >>
rect 1525 693 1554 722
<< m3 >>
rect 1525 693 1554 722
<< via2 >>
rect 1532 700 1547 715
<< m2 >>
rect 1101 1175 1131 1220
<< m3 >>
rect 1116 1160 1500 1190
<< m2 >>
rect 1485 864 1515 1175
<< m3 >>
rect 1500 849 1692 879
<< m2 >>
rect 1677 820 1707 864
<< m2 >>
rect 1109 1168 1138 1197
<< m3 >>
rect 1109 1168 1138 1197
<< via2 >>
rect 1116 1175 1131 1190
<< m2 >>
rect 1478 1153 1507 1182
<< m3 >>
rect 1478 1153 1507 1182
<< via2 >>
rect 1485 1160 1500 1175
<< m2 >>
rect 1493 857 1522 886
<< m3 >>
rect 1493 857 1522 886
<< via2 >>
rect 1500 864 1515 879
<< m2 >>
rect 1670 842 1699 871
<< m3 >>
rect 1670 842 1699 871
<< via2 >>
rect 1677 849 1692 864
<< m2 >>
rect 1869 740 1899 940
<< m3 >>
rect 1653 725 1884 755
<< m2 >>
rect 1638 673 1668 740
<< m3 >>
rect 1308 658 1653 688
<< m2 >>
rect 1293 540 1323 673
<< m2 >>
rect 1862 733 1891 762
<< m3 >>
rect 1862 733 1891 762
<< via2 >>
rect 1869 740 1884 755
<< m2 >>
rect 1646 718 1675 747
<< m3 >>
rect 1646 718 1675 747
<< via2 >>
rect 1653 725 1668 740
<< m2 >>
rect 1631 666 1660 695
<< m3 >>
rect 1631 666 1660 695
<< via2 >>
rect 1638 673 1653 688
<< m2 >>
rect 1301 651 1330 680
<< m3 >>
rect 1301 651 1330 680
<< via2 >>
rect 1308 658 1323 673
<< m2 >>
rect 1869 920 1899 940
<< m3 >>
rect 1860 905 1884 935
<< m2 >>
rect 1845 900 1875 920
<< m3 >>
rect 1740 885 1860 915
<< m2 >>
rect 1725 840 1755 900
<< m3 >>
rect 1692 825 1740 855
<< m2 >>
rect 1677 780 1707 840
<< m3 >>
rect 1668 765 1692 795
<< m2 >>
rect 1653 740 1683 780
<< m3 >>
rect 1596 725 1668 755
<< m2 >>
rect 1581 700 1611 740
<< m2 >>
rect 1862 913 1891 942
<< m3 >>
rect 1862 913 1891 942
<< via2 >>
rect 1869 920 1884 935
<< m2 >>
rect 1853 898 1882 927
<< m3 >>
rect 1853 898 1882 927
<< via2 >>
rect 1860 905 1875 920
<< m2 >>
rect 1838 893 1867 922
<< m3 >>
rect 1838 893 1867 922
<< via2 >>
rect 1845 900 1860 915
<< m2 >>
rect 1733 878 1762 907
<< m3 >>
rect 1733 878 1762 907
<< via2 >>
rect 1740 885 1755 900
<< m2 >>
rect 1718 833 1747 862
<< m3 >>
rect 1718 833 1747 862
<< via2 >>
rect 1725 840 1740 855
<< m2 >>
rect 1685 818 1714 847
<< m3 >>
rect 1685 818 1714 847
<< via2 >>
rect 1692 825 1707 840
<< m2 >>
rect 1670 773 1699 802
<< m3 >>
rect 1670 773 1699 802
<< via2 >>
rect 1677 780 1692 795
<< m2 >>
rect 1661 758 1690 787
<< m3 >>
rect 1661 758 1690 787
<< via2 >>
rect 1668 765 1683 780
<< m2 >>
rect 1646 733 1675 762
<< m3 >>
rect 1646 733 1675 762
<< via2 >>
rect 1653 740 1668 755
<< m2 >>
rect 1589 718 1618 747
<< m3 >>
rect 1589 718 1618 747
<< via2 >>
rect 1596 725 1611 740
<< m2 >>
rect 1005 2420 1035 2500
<< m3 >>
rect 1020 2405 1826 2435
<< m2 >>
rect 1811 2340 1841 2420
<< m3 >>
rect 1826 2325 1884 2355
<< m2 >>
rect 1013 2413 1042 2442
<< m3 >>
rect 1013 2413 1042 2442
<< via2 >>
rect 1020 2420 1035 2435
<< m2 >>
rect 1804 2398 1833 2427
<< m3 >>
rect 1804 2398 1833 2427
<< via2 >>
rect 1811 2405 1826 2420
<< m2 >>
rect 1819 2333 1848 2362
<< m3 >>
rect 1819 2333 1848 2362
<< via2 >>
rect 1826 2340 1841 2355
<< m3 >>
rect 1116 2605 1372 2635
<< m2 >>
rect 1357 2620 1387 2620
<< m3 >>
rect 1372 2605 1628 2635
<< m2 >>
rect 1613 2620 1643 2620
<< m3 >>
rect 1628 2605 1692 2635
<< m2 >>
rect 1101 2220 1131 2620
<< m3 >>
rect 1116 2605 1173 2635
<< m2 >>
rect 1158 2286 1188 2620
<< m3 >>
rect 1173 2271 1634 2301
<< m2 >>
rect 1619 2220 1649 2286
<< m3 >>
rect 1634 2205 1692 2235
<< m2 >>
rect 1151 2598 1180 2627
<< m3 >>
rect 1151 2598 1180 2627
<< via2 >>
rect 1158 2605 1173 2620
<< m2 >>
rect 1166 2279 1195 2308
<< m3 >>
rect 1166 2279 1195 2308
<< via2 >>
rect 1173 2286 1188 2301
<< m2 >>
rect 1612 2264 1641 2293
<< m3 >>
rect 1612 2264 1641 2293
<< via2 >>
rect 1619 2271 1634 2286
<< m2 >>
rect 1627 2213 1656 2242
<< m3 >>
rect 1627 2213 1656 2242
<< via2 >>
rect 1634 2220 1649 2235
<< m2 >>
rect 1677 2553 1707 2620
<< m3 >>
rect 1634 2538 1692 2568
<< m2 >>
rect 1619 2486 1649 2553
<< m3 >>
rect 1231 2471 1634 2501
<< m2 >>
rect 1216 2220 1246 2486
<< m3 >>
rect 1116 2205 1231 2235
<< m2 >>
rect 1670 2546 1699 2575
<< m3 >>
rect 1670 2546 1699 2575
<< via2 >>
rect 1677 2553 1692 2568
<< m2 >>
rect 1627 2531 1656 2560
<< m3 >>
rect 1627 2531 1656 2560
<< via2 >>
rect 1634 2538 1649 2553
<< m2 >>
rect 1612 2479 1641 2508
<< m3 >>
rect 1612 2479 1641 2508
<< via2 >>
rect 1619 2486 1634 2501
<< m2 >>
rect 1224 2464 1253 2493
<< m3 >>
rect 1224 2464 1253 2493
<< via2 >>
rect 1231 2471 1246 2486
<< m2 >>
rect 1209 2213 1238 2242
<< m3 >>
rect 1209 2213 1238 2242
<< via2 >>
rect 1216 2220 1231 2235
<< m2 >>
rect 1677 2620 1707 2620
<< m2 >>
rect 1677 2486 1707 2620
<< m2 >>
rect 1677 2486 1707 2486
<< m2 >>
rect 1677 2220 1707 2486
<< m3 >>
rect 1308 1925 1596 1955
<< m2 >>
rect 1581 1940 1611 2100
<< m2 >>
rect 1574 1933 1603 1962
<< m3 >>
rect 1574 1933 1603 1962
<< via2 >>
rect 1581 1940 1596 1955
<< m2 >>
rect 1101 2220 1131 2220
<< m3 >>
rect 1116 2205 1692 2235
<< m2 >>
rect 1677 2220 1707 2220
<< m3 >>
rect 1020 685 1164 715
<< m2 >>
rect 1149 638 1179 700
<< m3 >>
rect 1164 623 1308 653
<< m2 >>
rect 1293 601 1323 638
<< m3 >>
rect 1308 586 1596 616
<< m2 >>
rect 1581 589 1611 601
<< m3 >>
rect 1596 574 1644 604
<< m2 >>
rect 1629 576 1659 589
<< m3 >>
rect 1644 561 1788 591
<< m2 >>
rect 1773 540 1803 576
<< m3 >>
rect 1788 525 1884 555
<< m2 >>
rect 1142 678 1171 707
<< m3 >>
rect 1142 678 1171 707
<< via2 >>
rect 1149 685 1164 700
<< m2 >>
rect 1157 631 1186 660
<< m3 >>
rect 1157 631 1186 660
<< via2 >>
rect 1164 638 1179 653
<< m2 >>
rect 1286 616 1315 645
<< m3 >>
rect 1286 616 1315 645
<< via2 >>
rect 1293 623 1308 638
<< m2 >>
rect 1301 594 1330 623
<< m3 >>
rect 1301 594 1330 623
<< via2 >>
rect 1308 601 1323 616
<< m2 >>
rect 1574 582 1603 608
<< m3 >>
rect 1574 582 1603 608
<< via2 >>
rect 1581 589 1596 601
<< m2 >>
rect 1589 582 1618 608
<< m3 >>
rect 1589 582 1618 608
<< via2 >>
rect 1596 589 1611 601
<< m2 >>
rect 1622 569 1651 596
<< m3 >>
rect 1622 569 1651 596
<< via2 >>
rect 1629 576 1644 589
<< m2 >>
rect 1637 569 1666 596
<< m3 >>
rect 1637 569 1666 596
<< via2 >>
rect 1644 576 1659 589
<< m2 >>
rect 1766 554 1795 583
<< m3 >>
rect 1766 554 1795 583
<< via2 >>
rect 1773 561 1788 576
<< m2 >>
rect 1781 533 1810 562
<< m3 >>
rect 1781 533 1810 562
<< via2 >>
rect 1788 540 1803 555
<< labels >>
<< properties >>
<< end >>
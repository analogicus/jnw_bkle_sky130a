magic
tech sky130A
magscale 1 1
timestamp 1748204603
<< checkpaint >>
rect 0 0 1 1
use JNWATR_NCH_4C5F0  diff1_MN1 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 904
box 0 0 576 400
use JNWATR_NCH_4C5F0  diff1_MN2 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 904
box 0 0 576 400
use JNWATR_PCH_4C5F0  load1_MP5 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 3604
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP6 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 3204
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP  load1_MP6_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 3604
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP1 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  load1_MP1_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2164
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP2 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 2404
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT  load1_MP2_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 2164
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN4 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN4_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror2_MN3 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 504
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT  mirror2_MN3_TAPBOT ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 264
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN5 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 1304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN5_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 1704
box 0 0 576 240
use JNWATR_NCH_4C5F0  mirror1_MN6 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 1304
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP  mirror1_MN6_TAPTOP ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 1704
box 0 0 576 240
use JNWATR_PCH_4C5F0  load1_MP3 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 868 0 1 2804
box 0 0 576 400
use JNWATR_PCH_4C5F0  load1_MP4 ../JNW_ATR_SKY130A
timestamp 1748204603
transform 1 0 292 0 1 2804
box 0 0 576 400
<< m2 >>
rect 803 3225 1250 3255
<< m3 >>
rect 803 1321 833 3255
<< m2 >>
rect 674 1321 833 1351
<< m2 >>
rect 796 3218 840 3262
<< m3 >>
rect 796 3218 840 3262
<< via2 >>
rect 803 3225 833 3255
<< m2 >>
rect 796 1314 840 1358
<< m3 >>
rect 796 1314 840 1358
<< via2 >>
rect 803 1321 833 1351
<< m2 >>
rect 386 683 962 713
<< m2 >>
rect 244 2988 387 3018
<< m3 >>
rect 244 2588 274 3018
<< m2 >>
rect 244 2588 402 2618
<< m2 >>
rect 372 2588 978 2618
<< m2 >>
rect 948 2588 1266 2618
<< m3 >>
rect 1236 2588 1266 2858
<< m2 >>
rect 1236 2828 1410 2858
<< m3 >>
rect 1380 924 1410 2858
<< m2 >>
rect 1251 924 1410 954
<< m2 >>
rect 237 2981 281 3025
<< m3 >>
rect 237 2981 281 3025
<< via2 >>
rect 244 2988 274 3018
<< m2 >>
rect 237 2581 281 2625
<< m3 >>
rect 237 2581 281 2625
<< via2 >>
rect 244 2588 274 2618
<< m2 >>
rect 1229 2581 1273 2625
<< m3 >>
rect 1229 2581 1273 2625
<< via2 >>
rect 1236 2588 1266 2618
<< m2 >>
rect 1229 2821 1273 2865
<< m3 >>
rect 1229 2821 1273 2865
<< via2 >>
rect 1236 2828 1266 2858
<< m2 >>
rect 1373 2821 1417 2865
<< m3 >>
rect 1373 2821 1417 2865
<< via2 >>
rect 1380 2828 1410 2858
<< m2 >>
rect 1373 917 1417 961
<< m3 >>
rect 1373 917 1417 961
<< via2 >>
rect 1380 924 1410 954
<< m2 >>
rect 675 520 834 550
<< m3 >>
rect 804 520 834 1110
<< m2 >>
rect 596 1080 834 1110
<< m3 >>
rect 596 1080 626 1238
<< m2 >>
rect 468 1208 626 1238
<< m2 >>
rect 468 1208 1059 1238
<< m2 >>
rect 797 513 841 557
<< m3 >>
rect 797 513 841 557
<< via2 >>
rect 804 520 834 550
<< m2 >>
rect 797 1073 841 1117
<< m3 >>
rect 797 1073 841 1117
<< via2 >>
rect 804 1080 834 1110
<< m2 >>
rect 589 1073 633 1117
<< m3 >>
rect 589 1073 633 1117
<< via2 >>
rect 596 1080 626 1110
<< m2 >>
rect 589 1201 633 1245
<< m3 >>
rect 589 1201 633 1245
<< via2 >>
rect 596 1208 626 1238
<< m2 >>
rect 387 3388 978 3418
<< m2 >>
rect 948 3388 1410 3418
<< m3 >>
rect 1380 2988 1410 3418
<< m2 >>
rect 948 2988 1410 3018
<< m2 >>
rect 660 2988 978 3018
<< m3 >>
rect 660 2828 690 3018
<< m2 >>
rect 148 2828 690 2858
<< m3 >>
rect 148 924 178 2858
<< m2 >>
rect 148 924 675 954
<< m2 >>
rect 1373 3381 1417 3425
<< m3 >>
rect 1373 3381 1417 3425
<< via2 >>
rect 1380 3388 1410 3418
<< m2 >>
rect 1373 2981 1417 3025
<< m3 >>
rect 1373 2981 1417 3025
<< via2 >>
rect 1380 2988 1410 3018
<< m2 >>
rect 653 2981 697 3025
<< m3 >>
rect 653 2981 697 3025
<< via2 >>
rect 660 2988 690 3018
<< m2 >>
rect 653 2821 697 2865
<< m3 >>
rect 653 2821 697 2865
<< via2 >>
rect 660 2828 690 2858
<< m2 >>
rect 141 2821 185 2865
<< m3 >>
rect 141 2821 185 2865
<< via2 >>
rect 148 2828 178 2858
<< m2 >>
rect 141 917 185 961
<< m3 >>
rect 141 917 185 961
<< via2 >>
rect 148 924 178 954
<< m2 >>
rect 387 1484 978 1514
<< m2 >>
rect 660 1484 978 1514
<< m3 >>
rect 660 1484 690 2443
<< m2 >>
rect 653 1477 697 1521
<< m3 >>
rect 653 1477 697 1521
<< via2 >>
rect 660 1484 690 1514
<< locali >>
rect 100 3958 1636 4008
<< locali >>
rect 100 100 1636 150
<< m1 >>
rect 100 150 150 3958
<< m1 >>
rect 1586 150 1636 3958
<< locali >>
rect 93 3951 157 4015
<< m1 >>
rect 93 3951 157 4015
<< viali >>
rect 100 3958 150 4008
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1579 3951 1643 4015
<< m1 >>
rect 1579 3951 1643 4015
<< viali >>
rect 1586 3958 1636 4008
<< locali >>
rect 1579 93 1643 157
<< m1 >>
rect 1579 93 1643 157
<< viali >>
rect 1586 100 1636 150
<< locali >>
rect 0 4058 1736 4108
<< locali >>
rect 0 0 1736 50
<< m1 >>
rect 0 50 50 4058
<< m1 >>
rect 1686 50 1736 4058
<< locali >>
rect -7 4051 57 4115
<< m1 >>
rect -7 4051 57 4115
<< viali >>
rect 0 4058 50 4108
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1679 4051 1743 4115
<< m1 >>
rect 1679 4051 1743 4115
<< viali >>
rect 1686 4058 1736 4108
<< locali >>
rect 1679 -7 1743 57
<< m1 >>
rect 1679 -7 1743 57
<< viali >>
rect 1686 0 1736 50
<< locali >>
rect 244 3504 532 3544
<< locali >>
rect 628 3384 788 3424
<< locali >>
rect 820 3504 1108 3544
<< locali >>
rect 244 2704 532 2744
<< locali >>
rect 820 2704 1108 2744
<< locali >>
rect 1204 2584 1364 2624
<< locali >>
rect 244 804 532 844
<< locali >>
rect 820 804 1108 844
<< locali >>
rect 1204 684 1364 724
<< locali >>
rect 820 1604 1108 1644
<< locali >>
rect 1204 1484 1364 1524
<< locali >>
rect 244 1604 532 1644
<< locali >>
rect 820 3104 1108 3144
<< locali >>
rect 244 3104 532 3144
<< locali >>
rect 0 3676 1736 3772
<< locali >>
rect -7 3669 57 3779
<< m1 >>
rect -7 3669 57 3779
<< viali >>
rect 0 3676 50 3772
<< locali >>
rect 1679 3669 1743 3779
<< m1 >>
rect 1679 3669 1743 3779
<< viali >>
rect 1686 3676 1736 3772
<< locali >>
rect 0 2236 1736 2332
<< locali >>
rect -7 2229 57 2339
<< m1 >>
rect -7 2229 57 2339
<< viali >>
rect 0 2236 50 2332
<< locali >>
rect 1679 2229 1743 2339
<< m1 >>
rect 1679 2229 1743 2339
<< viali >>
rect 1686 2236 1736 2332
<< locali >>
rect 100 336 1636 432
<< locali >>
rect 93 329 157 439
<< m1 >>
rect 93 329 157 439
<< viali >>
rect 100 336 150 432
<< locali >>
rect 1579 329 1643 439
<< m1 >>
rect 1579 329 1643 439
<< viali >>
rect 1586 336 1636 432
<< locali >>
rect 100 1776 1636 1872
<< locali >>
rect 93 1769 157 1879
<< m1 >>
rect 93 1769 157 1879
<< viali >>
rect 100 1776 150 1872
<< locali >>
rect 1579 1769 1643 1879
<< m1 >>
rect 1579 1769 1643 1879
<< viali >>
rect 1586 1776 1636 1872
<< m1 >>
rect 1197 3217 1307 3271
<< m2 >>
rect 1197 3217 1307 3271
<< via1 >>
rect 1204 3224 1300 3264
<< m1 >>
rect 621 1317 731 1371
<< m2 >>
rect 621 1317 731 1371
<< via1 >>
rect 628 1324 724 1364
<< m1 >>
rect 365 677 411 731
<< m2 >>
rect 365 677 411 731
<< via1 >>
rect 372 684 404 724
<< m1 >>
rect 941 677 987 731
<< m2 >>
rect 941 677 987 731
<< via1 >>
rect 948 684 980 724
<< m1 >>
rect 1197 917 1307 971
<< m2 >>
rect 1197 917 1307 971
<< via1 >>
rect 1204 924 1300 964
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 365 2577 411 2631
<< m2 >>
rect 365 2577 411 2631
<< via1 >>
rect 372 2584 404 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 941 2577 987 2631
<< m2 >>
rect 941 2577 987 2631
<< via1 >>
rect 948 2584 980 2624
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< m3 >>
rect 1197 2817 1307 2871
<< via2 >>
rect 1204 2824 1300 2864
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 1197 2817 1307 2871
<< m2 >>
rect 1197 2817 1307 2871
<< via1 >>
rect 1204 2824 1300 2864
<< m1 >>
rect 365 2977 411 3031
<< m2 >>
rect 365 2977 411 3031
<< via1 >>
rect 372 2984 404 3024
<< m1 >>
rect 1005 1197 1115 1251
<< m2 >>
rect 1005 1197 1115 1251
<< via1 >>
rect 1012 1204 1108 1244
<< m1 >>
rect 429 1197 539 1251
<< m2 >>
rect 429 1197 539 1251
<< via1 >>
rect 436 1204 532 1244
<< m1 >>
rect 429 1197 539 1251
<< m2 >>
rect 429 1197 539 1251
<< via1 >>
rect 436 1204 532 1244
<< m1 >>
rect 621 517 731 571
<< m2 >>
rect 621 517 731 571
<< via1 >>
rect 628 524 724 564
<< m1 >>
rect 621 917 731 971
<< m2 >>
rect 621 917 731 971
<< via1 >>
rect 628 924 724 964
<< m1 >>
rect 365 3377 411 3431
<< m2 >>
rect 365 3377 411 3431
<< via1 >>
rect 372 3384 404 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 3377 987 3431
<< m2 >>
rect 941 3377 987 3431
<< via1 >>
rect 948 3384 980 3424
<< m1 >>
rect 941 2977 987 3031
<< m2 >>
rect 941 2977 987 3031
<< via1 >>
rect 948 2984 980 3024
<< m1 >>
rect 941 2977 987 3031
<< m2 >>
rect 941 2977 987 3031
<< via1 >>
rect 948 2984 980 3024
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< m3 >>
rect 621 2817 731 2871
<< via2 >>
rect 628 2824 724 2864
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2817 731 2871
<< m2 >>
rect 621 2817 731 2871
<< via1 >>
rect 628 2824 724 2864
<< m1 >>
rect 621 2417 731 2471
<< m2 >>
rect 621 2417 731 2471
<< m3 >>
rect 621 2417 731 2471
<< via2 >>
rect 628 2424 724 2464
<< via1 >>
rect 628 2424 724 2464
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 941 1477 987 1531
<< m2 >>
rect 941 1477 987 1531
<< via1 >>
rect 948 1484 980 1524
<< m1 >>
rect 365 1477 411 1531
<< m2 >>
rect 365 1477 411 1531
<< via1 >>
rect 372 1484 404 1524
use COMP2 U3_COMP2 
transform 1 0 1786 0 1 0
box 0 0 1786 4158
<< labels >>
flabel locali s 100 3958 1636 4008 0 FreeSans 400 0 0 0 VSS
port 42 nsew signal bidirectional
flabel locali s 0 4058 1736 4108 0 FreeSans 400 0 0 0 VDD
port 43 nsew signal bidirectional
flabel m1 s 948 1084 980 1124 0 FreeSans 400 0 0 0 VIP
port 44 nsew signal bidirectional
flabel m1 s 372 1084 404 1124 0 FreeSans 400 0 0 0 VIN
port 45 nsew signal bidirectional
flabel m2 s 803 3225 1250 3255 0 FreeSans 400 0 0 0 VO
port 46 nsew signal bidirectional
flabel m2 s 386 683 962 713 0 FreeSans 400 0 0 0 I_BIAS
port 47 nsew signal bidirectional
<< properties >>
<< end >>
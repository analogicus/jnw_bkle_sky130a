magic
tech sky130A
timestamp 1729602094
<< metal3 >>
rect 0 0 740 740
<< mimcap >>
rect 20 710 720 720
rect 20 30 30 710
rect 710 30 720 710
rect 20 20 720 30
<< mimcapcontact >>
rect 30 30 710 710
<< metal4 >>
rect 0 710 740 740
rect 0 30 30 710
rect 710 30 740 710
rect 0 0 740 30
<< labels >>
flabel metal4 s 0 0 740 50 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel metal3 s 0 0 740 50 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 740 740
<< end >>

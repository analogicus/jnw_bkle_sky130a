magic
tech sky130A
magscale 1 1
timestamp 1744591828
<< checkpaint >>
rect 0 0 0 0
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 1550
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP diff1_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 1950
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 806 0 1 1550
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP diff1_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 806 0 1 1950
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 550 0 1 2750
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 550 0 1 2510
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 2750
box 0 0 832 400
use JNWATR_PCH_12CTAPBOT load1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 2510
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 550 0 1 3550
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 550 0 1 3950
box 0 0 832 240
use JNWATR_PCH_12C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 3550
box 0 0 832 400
use JNWATR_PCH_12CTAPTOP load1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 3950
box 0 0 832 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 1150
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 806 0 1 1150
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 750
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror1_MN5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 510
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 806 0 1 750
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT mirror1_MN6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 806 0 1 510
box 0 0 576 240
use JNWATR_PCH_12C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 1382 0 1 3150
box 0 0 832 400
use JNWATR_PCH_12C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 550 0 1 3150
box 0 0 832 400
<< locali >>
rect 300 4300 2464 4400
<< locali >>
rect 300 300 2464 400
<< m1 >>
rect 300 400 400 4300
<< m1 >>
rect 2364 400 2464 4300
<< locali >>
rect 293 4293 407 4407
<< m1 >>
rect 293 4293 407 4407
<< viali >>
rect 300 4300 400 4400
<< locali >>
rect 293 293 407 407
<< m1 >>
rect 293 293 407 407
<< viali >>
rect 300 300 400 400
<< locali >>
rect 2357 4293 2471 4407
<< m1 >>
rect 2357 4293 2471 4407
<< viali >>
rect 2364 4300 2464 4400
<< locali >>
rect 2357 293 2471 407
<< m1 >>
rect 2357 293 2471 407
<< viali >>
rect 2364 300 2464 400
<< locali >>
rect 150 4450 2614 4550
<< locali >>
rect 150 150 2614 250
<< m1 >>
rect 150 250 250 4450
<< m1 >>
rect 2514 250 2614 4450
<< locali >>
rect 143 4443 257 4557
<< m1 >>
rect 143 4443 257 4557
<< viali >>
rect 150 4450 250 4550
<< locali >>
rect 143 143 257 257
<< m1 >>
rect 143 143 257 257
<< viali >>
rect 150 150 250 250
<< locali >>
rect 2507 4443 2621 4557
<< m1 >>
rect 2507 4443 2621 4557
<< viali >>
rect 2514 4450 2614 4550
<< locali >>
rect 2507 143 2621 257
<< m1 >>
rect 2507 143 2621 257
<< viali >>
rect 2514 150 2614 250
<< locali >>
rect 0 4600 2764 4700
<< locali >>
rect 0 0 2764 100
<< m1 >>
rect 0 100 100 4600
<< m1 >>
rect 2664 100 2764 4600
<< locali >>
rect -7 4593 107 4707
<< m1 >>
rect -7 4593 107 4707
<< viali >>
rect 0 4600 100 4700
<< locali >>
rect -7 -7 107 107
<< m1 >>
rect -7 -7 107 107
<< viali >>
rect 0 0 100 100
<< locali >>
rect 2657 4593 2771 4707
<< m1 >>
rect 2657 4593 2771 4707
<< viali >>
rect 2664 4600 2764 4700
<< locali >>
rect 2657 -7 2771 107
<< m1 >>
rect 2657 -7 2771 107
<< viali >>
rect 2664 0 2764 100
<< locali >>
rect 502 3050 790 3090
<< locali >>
rect 1142 2930 1302 2970
<< locali >>
rect 1334 3050 1622 3090
<< locali >>
rect 502 3850 790 3890
<< locali >>
rect 1334 3850 1622 3890
<< locali >>
rect 1974 3730 2134 3770
<< locali >>
rect 1334 1450 1622 1490
<< locali >>
rect 758 1450 1046 1490
<< locali >>
rect 1142 1330 1302 1370
<< locali >>
rect 1334 1050 1622 1090
<< locali >>
rect 1718 930 1878 970
<< locali >>
rect 758 1050 1046 1090
<< locali >>
rect 1334 3450 1622 3490
<< locali >>
rect 502 3450 790 3490
<< locali >>
rect 0 2022 2764 2118
<< locali >>
rect -7 2015 107 2125
<< m1 >>
rect -7 2015 107 2125
<< viali >>
rect 0 2022 100 2118
<< locali >>
rect 2657 2015 2771 2125
<< m1 >>
rect 2657 2015 2771 2125
<< viali >>
rect 2664 2022 2764 2118
<< locali >>
rect 150 2582 2614 2678
<< locali >>
rect 143 2575 257 2685
<< m1 >>
rect 143 2575 257 2685
<< viali >>
rect 150 2582 250 2678
<< locali >>
rect 2507 2575 2621 2685
<< m1 >>
rect 2507 2575 2621 2685
<< viali >>
rect 2514 2582 2614 2678
<< locali >>
rect 150 4022 2614 4118
<< locali >>
rect 143 4015 257 4125
<< m1 >>
rect 143 4015 257 4125
<< viali >>
rect 150 4022 250 4118
<< locali >>
rect 2507 4015 2621 4125
<< m1 >>
rect 2507 4015 2621 4125
<< viali >>
rect 2514 4022 2614 4118
<< locali >>
rect 0 582 2764 678
<< locali >>
rect -7 575 107 685
<< m1 >>
rect -7 575 107 685
<< viali >>
rect 0 582 100 678
<< locali >>
rect 2657 575 2771 685
<< m1 >>
rect 2657 575 2771 685
<< viali >>
rect 2664 582 2764 678
use COMP2 U2_COMP2 
transform 1 0 2814 0 1 0
box 0 0 2002 4450
use COMP2 U1_COMP2 
transform 1 0 4816 0 1 0
box 0 0 2002 4450
<< labels >>
flabel locali s 0 4600 2764 4700 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel locali s 150 4450 2614 4550 0 FreeSans 400 0 0 0 VDD
port 8 nsew signal bidirectional
<< properties >>
<< end >>
magic
tech sky130A
magscale 1 1
timestamp 1746029693
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 6440 4488 6490
<< locali >>
rect -100 -100 4488 -50
<< m1 >>
rect -100 -50 -50 6440
<< m1 >>
rect 4438 -50 4488 6440
<< locali >>
rect -107 6433 -43 6497
<< m1 >>
rect -107 6433 -43 6497
<< viali >>
rect -100 6440 -50 6490
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 4431 6433 4495 6497
<< m1 >>
rect 4431 6433 4495 6497
<< viali >>
rect 4438 6440 4488 6490
<< locali >>
rect 4431 -107 4495 -43
<< m1 >>
rect 4431 -107 4495 -43
<< viali >>
rect 4438 -100 4488 -50
<< locali >>
rect -200 6540 4588 6590
<< locali >>
rect -200 -200 4588 -150
<< m1 >>
rect -200 -150 -150 6540
<< m1 >>
rect 4538 -150 4588 6540
<< locali >>
rect -207 6533 -143 6597
<< m1 >>
rect -207 6533 -143 6597
<< viali >>
rect -200 6540 -150 6590
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 4531 6533 4595 6597
<< m1 >>
rect 4531 6533 4595 6597
<< viali >>
rect 4538 6540 4588 6590
<< locali >>
rect 4531 -207 4595 -143
<< m1 >>
rect 4531 -207 4595 -143
<< viali >>
rect 4538 -200 4588 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 4438 6440
<< labels >>
flabel locali s -100 6440 4488 6490 0 FreeSans 400 0 0 0 VDD
port 51 nsew signal bidirectional
flabel locali s -200 6540 4588 6590 0 FreeSans 400 0 0 0 VSS
port 52 nsew signal bidirectional
<< properties >>
<< end >>
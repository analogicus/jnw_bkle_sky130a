magic
tech sky130A
magscale 1 1
timestamp 1746183817
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP3<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<3>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP3<2>_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP3<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 1800
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP3<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 1800
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<3> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 2600
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<2> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 2600
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<1> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP4<0> ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 3400
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 3000
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 3400
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 776 0 1 -40
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 200 0 1 -40
box 0 0 576 240
use JNWTR_RPPO16 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1752 0 1 200
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1752 0 1 2020
box 0 0 2236 1720
use JNWTR_RPPO16 None_RH3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 1752 0 1 3795
box 0 0 2236 1720
use AALMISC_PNP_W3p40L3p40 None_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 4388 0 1 200
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 None_QP2 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 4388 0 1 990
box 0 0 670 670
<< m1 >>
rect 849 1573 895 1627
<< m2 >>
rect 849 1573 895 1627
<< via1 >>
rect 856 1580 888 1620
<< m1 >>
rect 273 1573 319 1627
<< m2 >>
rect 273 1573 319 1627
<< via1 >>
rect 280 1580 312 1620
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< m3 >>
rect 849 1973 895 2027
<< via2 >>
rect 856 1980 888 2020
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< via1 >>
rect 280 1980 312 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< m3 >>
rect 273 1973 319 2027
<< via2 >>
rect 280 1980 312 2020
<< via1 >>
rect 280 1980 312 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< via1 >>
rect 280 1980 312 2020
<< m1 >>
rect 273 2773 319 2827
<< m2 >>
rect 273 2773 319 2827
<< via1 >>
rect 280 2780 312 2820
<< m1 >>
rect 849 2773 895 2827
<< m2 >>
rect 849 2773 895 2827
<< via1 >>
rect 856 2780 888 2820
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< m3 >>
rect 849 2373 895 2427
<< via2 >>
rect 856 2380 888 2420
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< via1 >>
rect 280 2380 312 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< m3 >>
rect 273 2373 319 2427
<< via2 >>
rect 280 2380 312 2420
<< via1 >>
rect 280 2380 312 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< via1 >>
rect 280 2380 312 2420
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< m3 >>
rect 529 2613 639 2667
<< via2 >>
rect 536 2620 632 2660
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< m3 >>
rect 529 2613 639 2667
<< via2 >>
rect 536 2620 632 2660
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< m3 >>
rect 1105 2613 1215 2667
<< via2 >>
rect 1112 2620 1208 2660
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< m3 >>
rect 1105 2613 1215 2667
<< via2 >>
rect 1112 2620 1208 2660
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2213 1215 2267
<< m2 >>
rect 1105 2213 1215 2267
<< m3 >>
rect 1105 2213 1215 2267
<< via2 >>
rect 1112 2220 1208 2260
<< via1 >>
rect 1112 2220 1208 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< m3 >>
rect 529 2213 639 2267
<< via2 >>
rect 536 2220 632 2260
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< m3 >>
rect 529 2213 639 2267
<< via2 >>
rect 536 2220 632 2260
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 213 639 267
<< m2 >>
rect 529 213 639 267
<< via1 >>
rect 536 220 632 260
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< m3 >>
rect 1105 1413 1215 1467
<< via2 >>
rect 1112 1420 1208 1460
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< m3 >>
rect 1105 1413 1215 1467
<< via2 >>
rect 1112 1420 1208 1460
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< m3 >>
rect 1105 1413 1215 1467
<< via2 >>
rect 1112 1420 1208 1460
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 529 1413 639 1467
<< m2 >>
rect 529 1413 639 1467
<< m3 >>
rect 529 1413 639 1467
<< via2 >>
rect 536 1420 632 1460
<< via1 >>
rect 536 1420 632 1460
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< m3 >>
rect 1105 1813 1215 1867
<< via2 >>
rect 1112 1820 1208 1860
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< m3 >>
rect 1105 1813 1215 1867
<< via2 >>
rect 1112 1820 1208 1860
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< m3 >>
rect 529 1813 639 1867
<< via2 >>
rect 536 1820 632 1860
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< m3 >>
rect 529 1813 639 1867
<< via2 >>
rect 536 1820 632 1860
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< m3 >>
rect 849 373 895 427
<< via2 >>
rect 856 380 888 420
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< m3 >>
rect 849 373 895 427
<< via2 >>
rect 856 380 888 420
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< m3 >>
rect 1105 213 1215 267
<< via2 >>
rect 1112 220 1208 260
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< m3 >>
rect 1105 213 1215 267
<< via2 >>
rect 1112 220 1208 260
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 273 373 319 427
<< m2 >>
rect 273 373 319 427
<< via1 >>
rect 280 380 312 420
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< m3 >>
rect 913 1693 1023 1747
<< via2 >>
rect 920 1700 1016 1740
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< m3 >>
rect 337 1693 447 1747
<< via2 >>
rect 344 1700 440 1740
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< m3 >>
rect 913 2093 1023 2147
<< via2 >>
rect 920 2100 1016 2140
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 337 2093 447 2147
<< m2 >>
rect 337 2093 447 2147
<< via1 >>
rect 344 2100 440 2140
<< m1 >>
rect 337 2893 447 2947
<< m2 >>
rect 337 2893 447 2947
<< m3 >>
rect 337 2893 447 2947
<< via2 >>
rect 344 2900 440 2940
<< via1 >>
rect 344 2900 440 2940
<< m1 >>
rect 337 2893 447 2947
<< m2 >>
rect 337 2893 447 2947
<< via1 >>
rect 344 2900 440 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< m3 >>
rect 913 2893 1023 2947
<< via2 >>
rect 920 2900 1016 2940
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< m3 >>
rect 913 2493 1023 2547
<< via2 >>
rect 920 2500 1016 2540
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< m3 >>
rect 337 2493 447 2547
<< via2 >>
rect 344 2500 440 2540
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< m3 >>
rect 337 2493 447 2547
<< via2 >>
rect 344 2500 440 2540
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 529 3013 639 3067
<< m2 >>
rect 529 3013 639 3067
<< via1 >>
rect 536 3020 632 3060
<< m1 >>
rect 273 3173 319 3227
<< m2 >>
rect 273 3173 319 3227
<< via1 >>
rect 280 3180 312 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< m3 >>
rect 849 3173 895 3227
<< via2 >>
rect 856 3180 888 3220
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< m3 >>
rect 849 3173 895 3227
<< via2 >>
rect 856 3180 888 3220
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< via1 >>
rect 1112 3020 1208 3060
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< m3 >>
rect 1105 3013 1215 3067
<< via2 >>
rect 1112 3020 1208 3060
<< via1 >>
rect 1112 3020 1208 3060
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< via1 >>
rect 1112 3020 1208 3060
<< locali >>
rect 3655 1653 3813 1787
<< m1 >>
rect 3655 1653 3813 1787
<< m2 >>
rect 3655 1653 3813 1787
<< m3 >>
rect 3655 1653 3813 1787
<< via2 >>
rect 3662 1660 3806 1780
<< via1 >>
rect 3662 1660 3806 1780
<< viali >>
rect 3662 1660 3806 1780
<< locali >>
rect 1927 1653 2085 1787
<< m1 >>
rect 1927 1653 2085 1787
<< m2 >>
rect 1927 1653 2085 1787
<< m3 >>
rect 1927 1653 2085 1787
<< via2 >>
rect 1934 1660 2078 1780
<< via1 >>
rect 1934 1660 2078 1780
<< viali >>
rect 1934 1660 2078 1780
<< locali >>
rect 3655 3473 3813 3607
<< m1 >>
rect 3655 3473 3813 3607
<< m2 >>
rect 3655 3473 3813 3607
<< m3 >>
rect 3655 3473 3813 3607
<< via2 >>
rect 3662 3480 3806 3600
<< via1 >>
rect 3662 3480 3806 3600
<< viali >>
rect 3662 3480 3806 3600
<< locali >>
rect 1927 3473 2085 3607
<< m1 >>
rect 1927 3473 2085 3607
<< m2 >>
rect 1927 3473 2085 3607
<< m3 >>
rect 1927 3473 2085 3607
<< via2 >>
rect 1934 3480 2078 3600
<< via1 >>
rect 1934 3480 2078 3600
<< viali >>
rect 1934 3480 2078 3600
<< locali >>
rect 3655 5248 3813 5382
<< m1 >>
rect 3655 5248 3813 5382
<< m2 >>
rect 3655 5248 3813 5382
<< m3 >>
rect 3655 5248 3813 5382
<< via2 >>
rect 3662 5255 3806 5375
<< via1 >>
rect 3662 5255 3806 5375
<< viali >>
rect 3662 5255 3806 5375
<< m2 >>
rect 150 1582 293 1612
<< m3 >>
rect 150 1582 180 2012
<< m2 >>
rect 150 1982 308 2012
<< m3 >>
rect 278 1982 308 2012
<< m2 >>
rect 278 1982 884 2012
<< m3 >>
rect 854 1982 884 2012
<< m2 >>
rect 726 1982 884 2012
<< m3 >>
rect 726 1582 756 2012
<< m2 >>
rect 726 1582 869 1612
<< m1 >>
rect 849 1573 895 1627
<< m2 >>
rect 849 1573 895 1627
<< via1 >>
rect 856 1580 888 1620
<< m1 >>
rect 273 1573 319 1627
<< m2 >>
rect 273 1573 319 1627
<< via1 >>
rect 280 1580 312 1620
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 849 1973 895 2027
<< m2 >>
rect 849 1973 895 2027
<< via1 >>
rect 856 1980 888 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< via1 >>
rect 280 1980 312 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< via1 >>
rect 280 1980 312 2020
<< m1 >>
rect 273 1973 319 2027
<< m2 >>
rect 273 1973 319 2027
<< via1 >>
rect 280 1980 312 2020
<< m2 >>
rect 143 1575 187 1619
<< m3 >>
rect 143 1575 187 1619
<< via2 >>
rect 150 1582 180 1612
<< m2 >>
rect 143 1975 187 2019
<< m3 >>
rect 143 1975 187 2019
<< via2 >>
rect 150 1982 180 2012
<< m2 >>
rect 271 1975 315 2019
<< m3 >>
rect 271 1975 315 2019
<< via2 >>
rect 278 1982 308 2012
<< m2 >>
rect 271 1975 315 2019
<< m3 >>
rect 271 1975 315 2019
<< via2 >>
rect 278 1982 308 2012
<< m2 >>
rect 847 1975 891 2019
<< m3 >>
rect 847 1975 891 2019
<< via2 >>
rect 854 1982 884 2012
<< m2 >>
rect 847 1975 891 2019
<< m3 >>
rect 847 1975 891 2019
<< via2 >>
rect 854 1982 884 2012
<< m2 >>
rect 719 1975 763 2019
<< m3 >>
rect 719 1975 763 2019
<< via2 >>
rect 726 1982 756 2012
<< m2 >>
rect 719 1575 763 1619
<< m3 >>
rect 719 1575 763 1619
<< via2 >>
rect 726 1582 756 1612
<< m2 >>
rect 726 2782 869 2812
<< m3 >>
rect 726 2382 756 2812
<< m2 >>
rect 726 2382 884 2412
<< m3 >>
rect 854 2382 884 2412
<< m2 >>
rect 278 2382 884 2412
<< m3 >>
rect 278 2382 308 2412
<< m2 >>
rect 150 2382 308 2412
<< m3 >>
rect 150 2382 180 2812
<< m2 >>
rect 150 2782 293 2812
<< m1 >>
rect 273 2773 319 2827
<< m2 >>
rect 273 2773 319 2827
<< via1 >>
rect 280 2780 312 2820
<< m1 >>
rect 849 2773 895 2827
<< m2 >>
rect 849 2773 895 2827
<< via1 >>
rect 856 2780 888 2820
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 849 2373 895 2427
<< m2 >>
rect 849 2373 895 2427
<< via1 >>
rect 856 2380 888 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< via1 >>
rect 280 2380 312 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< via1 >>
rect 280 2380 312 2420
<< m1 >>
rect 273 2373 319 2427
<< m2 >>
rect 273 2373 319 2427
<< via1 >>
rect 280 2380 312 2420
<< m2 >>
rect 719 2775 763 2819
<< m3 >>
rect 719 2775 763 2819
<< via2 >>
rect 726 2782 756 2812
<< m2 >>
rect 719 2375 763 2419
<< m3 >>
rect 719 2375 763 2419
<< via2 >>
rect 726 2382 756 2412
<< m2 >>
rect 847 2375 891 2419
<< m3 >>
rect 847 2375 891 2419
<< via2 >>
rect 854 2382 884 2412
<< m2 >>
rect 847 2375 891 2419
<< m3 >>
rect 847 2375 891 2419
<< via2 >>
rect 854 2382 884 2412
<< m2 >>
rect 271 2375 315 2419
<< m3 >>
rect 271 2375 315 2419
<< via2 >>
rect 278 2382 308 2412
<< m2 >>
rect 271 2375 315 2419
<< m3 >>
rect 271 2375 315 2419
<< via2 >>
rect 278 2382 308 2412
<< m2 >>
rect 143 2375 187 2419
<< m3 >>
rect 143 2375 187 2419
<< via2 >>
rect 150 2382 180 2412
<< m2 >>
rect 143 2775 187 2819
<< m3 >>
rect 143 2775 187 2819
<< via2 >>
rect 150 2782 180 2812
<< m2 >>
rect 55 223 582 253
<< m3 >>
rect 55 223 85 2253
<< m2 >>
rect 55 2223 597 2253
<< m3 >>
rect 567 2223 597 2253
<< m3 >>
rect 567 2223 597 2653
<< m3 >>
rect 567 2623 597 2653
<< m2 >>
rect 567 2623 1173 2653
<< m3 >>
rect 1143 2623 1173 2653
<< m3 >>
rect 1143 2238 1173 2653
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 529 2613 639 2667
<< m2 >>
rect 529 2613 639 2667
<< via1 >>
rect 536 2620 632 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2613 1215 2667
<< m2 >>
rect 1105 2613 1215 2667
<< via1 >>
rect 1112 2620 1208 2660
<< m1 >>
rect 1105 2213 1215 2267
<< m2 >>
rect 1105 2213 1215 2267
<< via1 >>
rect 1112 2220 1208 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 2213 639 2267
<< m2 >>
rect 529 2213 639 2267
<< via1 >>
rect 536 2220 632 2260
<< m1 >>
rect 529 213 639 267
<< m2 >>
rect 529 213 639 267
<< via1 >>
rect 536 220 632 260
<< m2 >>
rect 48 216 92 260
<< m3 >>
rect 48 216 92 260
<< via2 >>
rect 55 223 85 253
<< m2 >>
rect 48 2216 92 2260
<< m3 >>
rect 48 2216 92 2260
<< via2 >>
rect 55 2223 85 2253
<< m2 >>
rect 560 2216 604 2260
<< m3 >>
rect 560 2216 604 2260
<< via2 >>
rect 567 2223 597 2253
<< m2 >>
rect 560 2616 604 2660
<< m3 >>
rect 560 2616 604 2660
<< via2 >>
rect 567 2623 597 2653
<< m2 >>
rect 1136 2616 1180 2660
<< m3 >>
rect 1136 2616 1180 2660
<< via2 >>
rect 1143 2623 1173 2653
<< m2 >>
rect 294 383 885 413
<< m3 >>
rect 855 383 885 413
<< m3 >>
rect 855 223 885 413
<< m2 >>
rect 855 223 1173 253
<< m3 >>
rect 1143 223 1173 253
<< m3 >>
rect 1143 223 1173 1453
<< m3 >>
rect 1143 1423 1173 1453
<< m3 >>
rect 1143 1423 1173 1853
<< m3 >>
rect 1143 1823 1173 1853
<< m2 >>
rect 567 1823 1173 1853
<< m3 >>
rect 567 1823 597 1853
<< m3 >>
rect 567 1438 597 1853
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 1105 1413 1215 1467
<< m2 >>
rect 1105 1413 1215 1467
<< via1 >>
rect 1112 1420 1208 1460
<< m1 >>
rect 529 1413 639 1467
<< m2 >>
rect 529 1413 639 1467
<< via1 >>
rect 536 1420 632 1460
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 1105 1813 1215 1867
<< m2 >>
rect 1105 1813 1215 1867
<< via1 >>
rect 1112 1820 1208 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 529 1813 639 1867
<< m2 >>
rect 529 1813 639 1867
<< via1 >>
rect 536 1820 632 1860
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 849 373 895 427
<< m2 >>
rect 849 373 895 427
<< via1 >>
rect 856 380 888 420
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 1105 213 1215 267
<< m2 >>
rect 1105 213 1215 267
<< via1 >>
rect 1112 220 1208 260
<< m1 >>
rect 273 373 319 427
<< m2 >>
rect 273 373 319 427
<< via1 >>
rect 280 380 312 420
<< m2 >>
rect 848 376 892 420
<< m3 >>
rect 848 376 892 420
<< via2 >>
rect 855 383 885 413
<< m2 >>
rect 848 216 892 260
<< m3 >>
rect 848 216 892 260
<< via2 >>
rect 855 223 885 253
<< m2 >>
rect 1136 216 1180 260
<< m3 >>
rect 1136 216 1180 260
<< via2 >>
rect 1143 223 1173 253
<< m2 >>
rect 1136 1816 1180 1860
<< m3 >>
rect 1136 1816 1180 1860
<< via2 >>
rect 1143 1823 1173 1853
<< m2 >>
rect 560 1816 604 1860
<< m3 >>
rect 560 1816 604 1860
<< via2 >>
rect 567 1823 597 1853
<< m2 >>
rect 392 3017 583 3047
<< m3 >>
rect 392 2537 422 3047
<< m2 >>
rect 376 2537 422 2567
<< m3 >>
rect 376 2505 406 2567
<< m2 >>
rect 408 2905 982 2935
<< m3 >>
rect 952 2905 982 2935
<< m2 >>
rect 952 2905 1318 2935
<< m3 >>
rect 1288 2505 1318 2935
<< m2 >>
rect 952 2505 1318 2535
<< m3 >>
rect 952 2505 982 2535
<< m2 >>
rect 952 2505 1318 2535
<< m3 >>
rect 1288 2105 1318 2535
<< m2 >>
rect 952 2105 1318 2135
<< m3 >>
rect 952 2105 982 2135
<< m2 >>
rect 952 2105 1318 2135
<< m3 >>
rect 1288 1705 1318 2135
<< m2 >>
rect 952 1705 1318 1735
<< m3 >>
rect 952 1705 982 1735
<< m2 >>
rect 376 1705 982 1735
<< m3 >>
rect 376 1705 406 1735
<< m2 >>
rect -40 1705 406 1735
<< m3 >>
rect -40 1705 -10 2135
<< m2 >>
rect -40 2105 391 2135
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 913 1693 1023 1747
<< m2 >>
rect 913 1693 1023 1747
<< via1 >>
rect 920 1700 1016 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 337 1693 447 1747
<< m2 >>
rect 337 1693 447 1747
<< via1 >>
rect 344 1700 440 1740
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 913 2093 1023 2147
<< m2 >>
rect 913 2093 1023 2147
<< via1 >>
rect 920 2100 1016 2140
<< m1 >>
rect 337 2093 447 2147
<< m2 >>
rect 337 2093 447 2147
<< via1 >>
rect 344 2100 440 2140
<< m1 >>
rect 337 2893 447 2947
<< m2 >>
rect 337 2893 447 2947
<< via1 >>
rect 344 2900 440 2940
<< m1 >>
rect 337 2893 447 2947
<< m2 >>
rect 337 2893 447 2947
<< via1 >>
rect 344 2900 440 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2893 1023 2947
<< m2 >>
rect 913 2893 1023 2947
<< via1 >>
rect 920 2900 1016 2940
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 913 2493 1023 2547
<< m2 >>
rect 913 2493 1023 2547
<< via1 >>
rect 920 2500 1016 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 337 2493 447 2547
<< m2 >>
rect 337 2493 447 2547
<< via1 >>
rect 344 2500 440 2540
<< m1 >>
rect 529 3013 639 3067
<< m2 >>
rect 529 3013 639 3067
<< via1 >>
rect 536 3020 632 3060
<< m2 >>
rect 385 3010 429 3054
<< m3 >>
rect 385 3010 429 3054
<< via2 >>
rect 392 3017 422 3047
<< m2 >>
rect 385 2530 429 2574
<< m3 >>
rect 385 2530 429 2574
<< via2 >>
rect 392 2537 422 2567
<< m2 >>
rect 369 2530 413 2574
<< m3 >>
rect 369 2530 413 2574
<< via2 >>
rect 376 2537 406 2567
<< m2 >>
rect 945 2898 989 2942
<< m3 >>
rect 945 2898 989 2942
<< via2 >>
rect 952 2905 982 2935
<< m2 >>
rect 945 2898 989 2942
<< m3 >>
rect 945 2898 989 2942
<< via2 >>
rect 952 2905 982 2935
<< m2 >>
rect 1281 2898 1325 2942
<< m3 >>
rect 1281 2898 1325 2942
<< via2 >>
rect 1288 2905 1318 2935
<< m2 >>
rect 1281 2498 1325 2542
<< m3 >>
rect 1281 2498 1325 2542
<< via2 >>
rect 1288 2505 1318 2535
<< m2 >>
rect 945 2498 989 2542
<< m3 >>
rect 945 2498 989 2542
<< via2 >>
rect 952 2505 982 2535
<< m2 >>
rect 945 2498 989 2542
<< m3 >>
rect 945 2498 989 2542
<< via2 >>
rect 952 2505 982 2535
<< m2 >>
rect 1281 2498 1325 2542
<< m3 >>
rect 1281 2498 1325 2542
<< via2 >>
rect 1288 2505 1318 2535
<< m2 >>
rect 1281 2098 1325 2142
<< m3 >>
rect 1281 2098 1325 2142
<< via2 >>
rect 1288 2105 1318 2135
<< m2 >>
rect 945 2098 989 2142
<< m3 >>
rect 945 2098 989 2142
<< via2 >>
rect 952 2105 982 2135
<< m2 >>
rect 945 2098 989 2142
<< m3 >>
rect 945 2098 989 2142
<< via2 >>
rect 952 2105 982 2135
<< m2 >>
rect 1281 2098 1325 2142
<< m3 >>
rect 1281 2098 1325 2142
<< via2 >>
rect 1288 2105 1318 2135
<< m2 >>
rect 1281 1698 1325 1742
<< m3 >>
rect 1281 1698 1325 1742
<< via2 >>
rect 1288 1705 1318 1735
<< m2 >>
rect 945 1698 989 1742
<< m3 >>
rect 945 1698 989 1742
<< via2 >>
rect 952 1705 982 1735
<< m2 >>
rect 945 1698 989 1742
<< m3 >>
rect 945 1698 989 1742
<< via2 >>
rect 952 1705 982 1735
<< m2 >>
rect 369 1698 413 1742
<< m3 >>
rect 369 1698 413 1742
<< via2 >>
rect 376 1705 406 1735
<< m2 >>
rect 369 1698 413 1742
<< m3 >>
rect 369 1698 413 1742
<< via2 >>
rect 376 1705 406 1735
<< m2 >>
rect -47 1698 -3 1742
<< m3 >>
rect -47 1698 -3 1742
<< via2 >>
rect -40 1705 -10 1735
<< m2 >>
rect -47 2098 -3 2142
<< m3 >>
rect -47 2098 -3 2142
<< via2 >>
rect -40 2105 -10 2135
<< m3 >>
rect 3717 1723 3747 3050
<< m2 >>
rect 1141 3020 3747 3050
<< m3 >>
rect 1141 3020 1171 3050
<< m2 >>
rect 853 3020 1171 3050
<< m3 >>
rect 853 3020 883 3210
<< m3 >>
rect 853 3180 883 3210
<< m2 >>
rect 292 3180 883 3210
<< m1 >>
rect 273 3173 319 3227
<< m2 >>
rect 273 3173 319 3227
<< via1 >>
rect 280 3180 312 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 849 3173 895 3227
<< m2 >>
rect 849 3173 895 3227
<< via1 >>
rect 856 3180 888 3220
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< via1 >>
rect 1112 3020 1208 3060
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< via1 >>
rect 1112 3020 1208 3060
<< m1 >>
rect 1105 3013 1215 3067
<< m2 >>
rect 1105 3013 1215 3067
<< via1 >>
rect 1112 3020 1208 3060
<< locali >>
rect 3655 1653 3813 1787
<< m1 >>
rect 3655 1653 3813 1787
<< viali >>
rect 3662 1660 3806 1780
<< m2 >>
rect 3710 3013 3754 3057
<< m3 >>
rect 3710 3013 3754 3057
<< via2 >>
rect 3717 3020 3747 3050
<< m2 >>
rect 1134 3013 1178 3057
<< m3 >>
rect 1134 3013 1178 3057
<< via2 >>
rect 1141 3020 1171 3050
<< m2 >>
rect 1134 3013 1178 3057
<< m3 >>
rect 1134 3013 1178 3057
<< via2 >>
rect 1141 3020 1171 3050
<< m2 >>
rect 846 3013 890 3057
<< m3 >>
rect 846 3013 890 3057
<< via2 >>
rect 853 3020 883 3050
<< m2 >>
rect 846 3173 890 3217
<< m3 >>
rect 846 3173 890 3217
<< via2 >>
rect 853 3180 883 3210
<< m3 >>
rect 1986 1718 2016 3349
<< m2 >>
rect 1986 3319 3744 3349
<< m3 >>
rect 3714 3319 3744 3542
<< locali >>
rect 1927 1653 2085 1787
<< m1 >>
rect 1927 1653 2085 1787
<< viali >>
rect 1934 1660 2078 1780
<< locali >>
rect 3655 3473 3813 3607
<< m1 >>
rect 3655 3473 3813 3607
<< viali >>
rect 3662 3480 3806 3600
<< m2 >>
rect 1979 3312 2023 3356
<< m3 >>
rect 1979 3312 2023 3356
<< via2 >>
rect 1986 3319 2016 3349
<< m2 >>
rect 3707 3312 3751 3356
<< m3 >>
rect 3707 3312 3751 3356
<< via2 >>
rect 3714 3319 3744 3349
<< m3 >>
rect 1986 3540 2016 4483
<< m2 >>
rect 1986 4453 3744 4483
<< m3 >>
rect 3714 4453 3744 5300
<< locali >>
rect 1927 3473 2085 3607
<< m1 >>
rect 1927 3473 2085 3607
<< viali >>
rect 1934 3480 2078 3600
<< locali >>
rect 3655 5248 3813 5382
<< m1 >>
rect 3655 5248 3813 5382
<< viali >>
rect 3662 5255 3806 5375
<< m2 >>
rect 1979 4446 2023 4490
<< m3 >>
rect 1979 4446 2023 4490
<< via2 >>
rect 1986 4453 2016 4483
<< m2 >>
rect 3707 4446 3751 4490
<< m3 >>
rect 3707 4446 3751 4490
<< via2 >>
rect 3714 4453 3744 4483
<< locali >>
rect 100 5565 5158 5615
<< locali >>
rect 100 100 5158 150
<< m1 >>
rect 100 150 150 5565
<< m1 >>
rect 5108 150 5158 5565
<< locali >>
rect 93 5558 157 5622
<< m1 >>
rect 93 5558 157 5622
<< viali >>
rect 100 5565 150 5615
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 5101 5558 5165 5622
<< m1 >>
rect 5101 5558 5165 5622
<< viali >>
rect 5108 5565 5158 5615
<< locali >>
rect 5101 93 5165 157
<< m1 >>
rect 5101 93 5165 157
<< viali >>
rect 5108 100 5158 150
<< locali >>
rect 0 5665 5258 5715
<< locali >>
rect 0 0 5258 50
<< m1 >>
rect 0 50 50 5665
<< m1 >>
rect 5208 50 5258 5665
<< locali >>
rect -7 5658 57 5722
<< m1 >>
rect -7 5658 57 5722
<< viali >>
rect 0 5665 50 5715
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 5201 5658 5265 5722
<< m1 >>
rect 5201 5658 5265 5722
<< viali >>
rect 5208 5665 5258 5715
<< locali >>
rect 5201 -7 5265 57
<< m1 >>
rect 5201 -7 5265 57
<< viali >>
rect 5208 0 5258 50
<< locali >>
rect 152 3300 440 3340
<< locali >>
rect 728 3300 1016 3340
<< locali >>
rect 1112 3180 1272 3220
<< locali >>
rect 728 500 1016 540
<< locali >>
rect 1112 380 1272 420
<< locali >>
rect 152 500 440 540
<< locali >>
rect 100 1232 1352 1328
<< locali >>
rect 93 1225 157 1335
<< m1 >>
rect 93 1225 157 1335
<< viali >>
rect 100 1232 150 1328
<< locali >>
rect 100 3472 1352 3568
<< locali >>
rect 93 3465 157 3575
<< m1 >>
rect 93 3465 157 3575
<< viali >>
rect 100 3472 150 3568
<< locali >>
rect 0 672 1352 768
<< locali >>
rect -7 665 57 775
<< m1 >>
rect -7 665 57 775
<< viali >>
rect 0 672 50 768
<< locali >>
rect 0 32 1352 128
<< locali >>
rect -7 25 57 135
<< m1 >>
rect -7 25 57 135
<< viali >>
rect 0 32 50 128
<< locali >>
rect 1760 5255 2078 5375
<< locali >>
rect 1552 1864 4188 1920
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 1857 1609 1927
<< m1 >>
rect 1545 1857 1609 1927
<< viali >>
rect 1552 1864 1602 1920
<< locali >>
rect 4131 1857 4195 1927
<< m1 >>
rect 4131 1857 4195 1927
<< viali >>
rect 4138 1864 4188 1920
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 1857 1609 1927
<< m1 >>
rect 1545 1857 1609 1927
<< viali >>
rect 1552 1864 1602 1920
<< locali >>
rect 1552 200 4188 256
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 193 1609 263
<< m1 >>
rect 1545 193 1609 263
<< viali >>
rect 1552 200 1602 256
<< locali >>
rect 4131 193 4195 263
<< m1 >>
rect 4131 193 4195 263
<< viali >>
rect 4138 200 4188 256
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 193 1609 263
<< m1 >>
rect 1545 193 1609 263
<< viali >>
rect 1552 200 1602 256
<< locali >>
rect 1552 3684 4188 3740
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 3677 1609 3747
<< m1 >>
rect 1545 3677 1609 3747
<< viali >>
rect 1552 3684 1602 3740
<< locali >>
rect 4131 3677 4195 3747
<< m1 >>
rect 4131 3677 4195 3747
<< viali >>
rect 4138 3684 4188 3740
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 3677 1609 3747
<< m1 >>
rect 1545 3677 1609 3747
<< viali >>
rect 1552 3684 1602 3740
<< locali >>
rect 1552 2020 4188 2076
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 2013 1609 2083
<< m1 >>
rect 1545 2013 1609 2083
<< viali >>
rect 1552 2020 1602 2076
<< locali >>
rect 4131 2013 4195 2083
<< m1 >>
rect 4131 2013 4195 2083
<< viali >>
rect 4138 2020 4188 2076
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 2013 1609 2083
<< m1 >>
rect 1545 2013 1609 2083
<< viali >>
rect 1552 2020 1602 2076
<< locali >>
rect 1552 5459 4188 5515
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 5452 1609 5522
<< m1 >>
rect 1545 5452 1609 5522
<< viali >>
rect 1552 5459 1602 5515
<< locali >>
rect 4131 5452 4195 5522
<< m1 >>
rect 4131 5452 4195 5522
<< viali >>
rect 4138 5459 4188 5515
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 5452 1609 5522
<< m1 >>
rect 1545 5452 1609 5522
<< viali >>
rect 1552 5459 1602 5515
<< locali >>
rect 1552 3795 4188 3851
<< m1 >>
rect 1552 0 1602 5715
<< m1 >>
rect 4138 0 4188 5715
<< locali >>
rect 1545 3788 1609 3858
<< m1 >>
rect 1545 3788 1609 3858
<< viali >>
rect 1552 3795 1602 3851
<< locali >>
rect 4131 3788 4195 3858
<< m1 >>
rect 4131 3788 4195 3858
<< viali >>
rect 4138 3795 4188 3851
<< locali >>
rect 4131 -7 4195 57
<< m1 >>
rect 4131 -7 4195 57
<< viali >>
rect 4138 0 4188 50
<< locali >>
rect 4131 5658 4195 5722
<< m1 >>
rect 4131 5658 4195 5722
<< viali >>
rect 4138 5665 4188 5715
<< locali >>
rect 1545 -7 1609 57
<< m1 >>
rect 1545 -7 1609 57
<< viali >>
rect 1552 0 1602 50
<< locali >>
rect 1545 5658 1609 5722
<< m1 >>
rect 1545 5658 1609 5722
<< viali >>
rect 1552 5665 1602 5715
<< locali >>
rect 1545 3788 1609 3858
<< m1 >>
rect 1545 3788 1609 3858
<< viali >>
rect 1552 3795 1602 3851
<< locali >>
rect 4388 846 5258 870
<< locali >>
rect 5201 839 5265 877
<< m1 >>
rect 5201 839 5265 877
<< viali >>
rect 5208 846 5258 870
<< locali >>
rect 4388 200 5258 224
<< locali >>
rect 5201 193 5265 231
<< m1 >>
rect 5201 193 5265 231
<< viali >>
rect 5208 200 5258 224
<< locali >>
rect 4388 1636 5258 1660
<< locali >>
rect 5201 1629 5265 1667
<< m1 >>
rect 5201 1629 5265 1667
<< viali >>
rect 5208 1636 5258 1660
<< locali >>
rect 4388 990 5258 1014
<< locali >>
rect 5201 983 5265 1021
<< m1 >>
rect 5201 983 5265 1021
<< viali >>
rect 5208 990 5258 1014
<< labels >>
flabel m2 s 150 1582 293 1612 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel m2 s 726 2782 869 2812 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel locali s 100 5565 5158 5615 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel locali s 0 5665 5258 5715 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel m2 s 55 223 582 253 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>
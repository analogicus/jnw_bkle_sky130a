magic
tech sky130A
magscale 1 1
timestamp 1745853979
<< checkpaint >>
rect 0 0 1 1
<< locali >>
rect -100 10040 2936 10090
<< locali >>
rect -100 -100 2936 -50
<< m1 >>
rect -100 -50 -50 10040
<< m1 >>
rect 2886 -50 2936 10040
<< locali >>
rect -107 10033 -43 10097
<< m1 >>
rect -107 10033 -43 10097
<< viali >>
rect -100 10040 -50 10090
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 2879 10033 2943 10097
<< m1 >>
rect 2879 10033 2943 10097
<< viali >>
rect 2886 10040 2936 10090
<< locali >>
rect 2879 -107 2943 -43
<< m1 >>
rect 2879 -107 2943 -43
<< viali >>
rect 2886 -100 2936 -50
<< locali >>
rect -200 10140 3036 10190
<< locali >>
rect -200 -200 3036 -150
<< m1 >>
rect -200 -150 -150 10140
<< m1 >>
rect 2986 -150 3036 10140
<< locali >>
rect -207 10133 -143 10197
<< m1 >>
rect -207 10133 -143 10197
<< viali >>
rect -200 10140 -150 10190
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 2979 10133 3043 10197
<< m1 >>
rect 2979 10133 3043 10197
<< viali >>
rect 2986 10140 3036 10190
<< locali >>
rect 2979 -207 3043 -143
<< m1 >>
rect 2979 -207 3043 -143
<< viali >>
rect 2986 -200 3036 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 2886 10040
<< labels >>
flabel locali s -100 10040 2936 10090 0 FreeSans 400 0 0 0 VDD
port 51 nsew signal bidirectional
flabel locali s -200 10140 3036 10190 0 FreeSans 400 0 0 0 VSS
port 52 nsew signal bidirectional
<< properties >>
<< end >>                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< m3 >>
rect 629 7503 739 7557
<< via2 >>
rect 636 7510 732 7550
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< m3 >>
rect 629 7503 739 7557
<< via2 >>
rect 636 7510 732 7550
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< m3 >>
rect 629 6303 739 6357
<< via2 >>
rect 636 6310 732 6350
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< m3 >>
rect 629 6303 739 6357
<< via2 >>
rect 636 6310 732 6350
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 949 6463 995 6517
<< m2 >>
rect 949 6463 995 6517
<< m3 >>
rect 949 6463 995 6517
<< via2 >>
rect 956 6470 988 6510
<< via1 >>
rect 956 6470 988 6510
<< m1 >>
rect 373 9263 419 9317
<< m2 >>
rect 373 9263 419 9317
<< via1 >>
rect 380 9270 412 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< m3 >>
rect 949 9263 995 9317
<< via2 >>
rect 956 9270 988 9310
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< m3 >>
rect 949 9263 995 9317
<< via2 >>
rect 956 9270 988 9310
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 949 9263 995 9317
<< m2 >>
rect 949 9263 995 9317
<< via1 >>
rect 956 9270 988 9310
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< m3 >>
rect 1205 9103 1315 9157
<< via2 >>
rect 1212 9110 1308 9150
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< m3 >>
rect 1205 9103 1315 9157
<< via2 >>
rect 1212 9110 1308 9150
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< locali >>
rect 2203 1953 2361 2087
<< m1 >>
rect 2203 1953 2361 2087
<< m2 >>
rect 2203 1953 2361 2087
<< via1 >>
rect 2210 1960 2354 2080
<< viali >>
rect 2210 1960 2354 2080
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< m2 >>
rect 475 1953 633 2087
<< m3 >>
rect 475 1953 633 2087
<< via2 >>
rect 482 1960 626 2080
<< via1 >>
rect 482 1960 626 2080
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< m2 >>
rect 2203 3773 2361 3907
<< via1 >>
rect 2210 3780 2354 3900
<< viali >>
rect 2210 3780 2354 3900
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< m2 >>
rect 475 3773 633 3907
<< m3 >>
rect 475 3773 633 3907
<< via2 >>
rect 482 3780 626 3900
<< via1 >>
rect 482 3780 626 3900
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< m2 >>
rect 2203 5623 2361 5757
<< m3 >>
rect 2203 5623 2361 5757
<< via2 >>
rect 2210 5630 2354 5750
<< via1 >>
rect 2210 5630 2354 5750
<< viali >>
rect 2210 5630 2354 5750
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< m3 >>
rect 1013 8183 1123 8237
<< via2 >>
rect 1020 8190 1116 8230
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< m3 >>
rect 1013 8183 1123 8237
<< via2 >>
rect 1020 8190 1116 8230
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< m3 >>
rect 437 7783 547 7837
<< via2 >>
rect 444 7790 540 7830
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 10205 8703 1315 8757
<< m3 >>
rect 1205 8703 1315 8757
<< via2 >>
rect 1212 8710 1308 8750
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 1205 8703 1315 8757
<< m2 >>
rect 1205 8703 1315 8757
<< m3 >>
rect 1205 8703 1315 8757
<< via2 >>
rect 1212 8710 1308 8750
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 1205 8703 1315 8757
<< m2 >>
rect 1205 8703 1315 8757
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 629 8703 739 8757
<< m2 >>
rect 629 8703 739 8757
<< m3 >>
rect 629 8703 739 8757
<< via2 >>
rect 636 8710 732 8750
<< via1 >>
rect 636 8710 732 8750
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< m3 >>
rect 1205 6303 1315 6357
<< via2 >>
rect 1212 6310 1308 6350
<< via1 >>
rect 1212 6310 1308 6350
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< m2 >>
rect 475 1953 633 2087
<< m3 >>
rect 475 1953 633 2087
<< via2 >>
rect 482 1960 626 2080
<< via1 >>
rect 482 1960 626 2080
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< m2 >>
rect 2203 3773 2361 3907
<< via1 >>
rect 2210 3780 2354 3900
<< viali >>
rect 2210 3780 2354 3900
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< m2 >>
rect 475 3773 633 3907
<< m3 >>
rect 475 3773 633 3907
<< via2 >>
rect 482 3780 626 3900
<< via1 >>
rect 482 3780 626 3900
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< m2 >>
rect 2203 5623 2361 5757
<< via1 >>
rect 2210 5630 2354 5750
<< viali >>
rect 2210 5630 2354 5750
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< m3 >>
rect 1013 7783 1123 7837
<< via2 >>
rect 1020 7790 1116 7830
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< m3 >>
rect 1013 7783 1123 7837
<< via2 >>
rect 1020 7790 1116 7830
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< m3 >>
rect 437 8183 547 8237
<< via2 >>
rect 444 8190 540 8230
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< m3 >>
rect 437 8183 547 8237
<< via2 >>
rect 444 8190 540 8230
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 1013 8583 1123 8637
<< m2 >>
rect 1013 8583 1123 8637
<< via1 >>
rect 1020 8590 1116 8630
<< m1 >>
rect 437 8583 547 8637
<< m2 >>
rect 437 8583 547 8637
<< m3 >>
rect 437 8583 547 8637
<< via2 >>
rect 444 8590 540 8630
<< via1 >>
rect 444 8590 540 8630
<< m1 >>
rect 437 8583 547 8637
<< m2 >>
rect 437 8583 547 8637
<< via1 >>
rect 444 8590 540 8630
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< m3 >>
rect 1013 8983 1123 9037
<< via2 >>
rect 1020 8990 1116 9030
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 437 8983 547 9037
<< m2 >>
rect 437 8983 547 9037
<< via1 >>
rect 444 8990 540 9030
<< m1 >>
rect 437 8983 547 9037
<< m2 >>
rect 437 8983 547 9037
<< m3 >>
rect 437 8983 547 9037
<< via2 >>
rect 444 8990 540 9030
<< via1 >>
rect 444 8990 540 9030
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< m3 >>
rect 1205 9103 1315 9157
<< via2 >>
rect 1212 9110 1308 9150
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m3 >>
rect 955 6313 985 6488
<< m2 >>
rect 667 6313 985 6343
<< m3 >>
rect 667 6313 697 6343
<< m3 >>
rect 667 6313 697 7543
<< m3 >>
rect 667 7513 697 7543
<< m2 >>
rect 667 7513 841 7543
<< m3 >>
rect 811 7513 841 7703
<< m2 >>
rect 667 7673 841 7703
<< m3 >>
rect 667 7673 697 7943
<< m3 >>
rect 667 7913 697 7943
<< m2 >>
rect 667 7913 1273 7943
<< m3 >>
rect 1243 7913 1273 7943
<< m3 >>
rect 1243 7528 1273 7943
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 629 7503 739 7557
<< m2 >>
rect 629 7503 739 7557
<< via1 >>
rect 636 7510 732 7550
<< m1 >>
rect 1205 7503 1315 7557
<< m2 >>
rect 1205 7503 1315 7557
<< via1 >>
rect 1212 7510 1308 7550
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 1205 7903 1315 7957
<< m2 >>
rect 1205 7903 1315 7957
<< via1 >>
rect 1212 7910 1308 7950
<< m1 >>
rect 629 7903 739 7957
<< m2 >>
rect 629 7903 739 7957
<< via1 >>
rect 636 7910 732 7950
<< m1 >>
rect 629 7903 739 7957
<< m2 >>
rect 629 7903 739 7957
<< via1 >>
rect 636 7910 732 7950
<< m1 >>
rect 629 7903 739 7957
<< m2 >>
rect 629 7903 739 7957
<< via1 >>
rect 636 7910 732 7950
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 629 6303 739 6357
<< m2 >>
rect 629 6303 739 6357
<< via1 >>
rect 636 6310 732 6350
<< m1 >>
rect 949 6463 995 6517
<< m2 >>
rect 949 6463 995 6517
<< via1 >>
rect 956 6470 988 6510
<< m2 >>
rect 948 6306 992 6350
<< m3 >>
rect 948 6306 992 6350
<< via2 >>
rect 955 6313 985 6343
<< m2 >>
rect 660 6306 704 6350
<< m3 >>
rect 660 6306 704 6350
<< via2 >>
rect 667 6313 697 6343
<< m2 >>
rect 660 7506 704 7550
<< m3 >>
rect 660 7506 704 7550
<< via2 >>
rect 667 7513 697 7543
<< m2 >>
rect 804 7506 848 7550
<< m3 >>
rect 804 7506 848 7550
<< via2 >>
rect 811 7513 841 7543
<< m2 >>
rect 804 7666 848 7710
<< m3 >>
rect 804 7666 848 7710
<< via2 >>
rect 811 7673 841 7703
<< m2 >>
rect 660 7666 704 7710
<< m3 >>
rect 660 7666 704 7710
<< via2 >>
rect 667 7673 697 7703
<< m2 >>
rect 660 7906 704 7950
<< m3 >>
rect 660 7906 704 7950
<< via2 >>
rect 667 7913 697 7943
<< m2 >>
rect 1236 7906 1280 7950
<< m3 >>
rect 1236 7906 1280 7950
<< via2 >>
rect 1243 7913 1273 7943
<< m2 >>
rect 234 8473 393 8503
<< m3 >>
rect 234 8473 264 8759
<< m2 >>
rect 234 8729 408 8759
<< m3 >>
rect 378 8729 408 8903
<< m3 >>
rect 378 8873 408 8903
<< m2 >>
rect 378 8873 984 8903
<< m3 >>
rect 954 8873 984 8903
<< m3 >>
rect 954 8713 984 8903
<< m2 >>
rect 810 8713 984 8743
<< m3 >>
rect 810 8473 840 8743
<< m2 >>
rect 810 8473 969 8503
<< m1 >>
rect 949 8463 995 8517
<< m2 >>
rect 949 8463 995 8517
<< via1 >>
rect 956 8470 988 8510
<< m1 >>
rect 373 8463 419 8517
<< m2 >>
rect 373 8463 419 8517
<< via1 >>
rect 380 8470 412 8510
<< m1 >>
rect 949 8863 995 8917
<< m2 >>
rect 949 8863 995 8917
<< via1 >>
rect 956 8870 988 8910
<< m1 >>
rect 949 8863 995 8917
<< m2 >>
rect 949 8863 995 8917
<< via1 >>
rect 956 8870 988 8910
<< m1 >>
rect 949 8863 995 8917
<< m2 >>
rect 949 8863 995 8917
<< via1 >>
rect 956 8870 988 8910
<< m1 >>
rect 373 8863 419 8917
<< m2 >>
rect 373 8863 419 8917
<< via1 >>
rect 380 8870 412 8910
<< m1 >>
rect 373 8863 419 8917
<< m2 >>
rect 373 8863 419 8917
<< via1 >>
rect 380 8870 412 8910
<< m1 >>
rect 373 8863 419 8917
<< m2 >>
rect 373 8863 419 8917
<< via1 >>
rect 380 8870 412 8910
<< m2 >>
rect 227 8466 271 8510
<< m3 >>
rect 227 8466 271 8510
<< via2 >>
rect 234 8473 264 8503
<< m2 >>
rect 227 8722 271 8766
<< m3 >>
rect 227 8722 271 8766
<< via2 >>
rect 234 8729 264 8759
<< m2 >>
rect 371 8722 415 8766
<< m3 >>
rect 371 8722 415 8766
<< via2 >>
rect 378 8729 408 8759
<< m2 >>
rect 371 8866 415 8910
<< m3 >>
rect 371 8866 415 8910
<< via2 >>
rect 378 8873 408 8903
<< m2 >>
rect 947 8866 991 8910
<< m3 >>
rect 947 8866 991 8910
<< via2 >>
rect 954 8873 984 8903
<< m2 >>
rect 947 8706 991 8750
<< m3 >>
rect 947 8706 991 8750
<< via2 >>
rect 954 8713 984 8743
<< m2 >>
rect 803 8706 847 8750
<< m3 >>
rect 803 8706 847 8750
<< via2 >>
rect 810 8713 840 8743
<< m2 >>
rect 803 8466 847 8510
<< m3 >>
rect 803 8466 847 8510
<< via2 >>
rect 810 8473 840 8503
<< m2 >>
rect 969 7673 1416 7703
<< m3 >>
rect 1386 7673 1416 8103
<< m2 >>
rect 954 8073 1416 8103
<< m3 >>
rect 954 7673 984 8103
<< m3 >>
rect 954 7401 984 7703
<< m2 >>
rect 442 7401 984 7431
<< m3 >>
rect 442 7401 472 7799
<< m2 >>
rect 234 7769 472 7799
<< m3 >>
rect 234 7769 264 7943
<< m2 >>
rect 234 7913 408 7943
<< m3 >>
rect 378 7913 408 8103
<< m3 >>
rect 378 8073 408 8103
<< m3 >>
rect 378 7913 408 8103
<< m2 >>
rect 234 7913 408 7943
<< m3 >>
rect 234 7673 264 7943
<< m2 >>
rect 234 7673 393 7703
<< m1 >>
rect 373 7663 419 7717
<< m2 >>
rect 373 7663 419 7717
<< via1 >>
rect 380 7670 412 7710
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 437 7783 547 7837
<< m2 >>
rect 437 7783 547 7837
<< via1 >>
rect 444 7790 540 7830
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 7663 995 7717
<< m2 >>
rect 949 7663 995 7717
<< via1 >>
rect 956 7670 988 7710
<< m1 >>
rect 949 8063 995 8117
<< m2 >>
rect 949 8063 995 8117
<< via1 >>
rect 956 8070 988 8110
<< m1 >>
rect 949 8063 995 8117
<< m2 >>
rect 949 8063 995 8117
<< via1 >>
rect 956 8070 988 8110
<< m1 >>
rect 373 8063 419 8117
<< m2 >>
rect 373 8063 419 8117
<< via1 >>
rect 380 8070 412 8110
<< m1 >>
rect 373 8063 419 8117
<< m2 >>
rect 373 8063 419 8117
<< via1 >>
rect 380 8070 412 8110
<< m1 >>
rect 373 8063 419 8117
<< m2 >>
rect 373 8063 419 8117
<< via1 >>
rect 380 8070 412 8110
<< m2 >>
rect 1379 7666 1423 7710
<< m3 >>
rect 1379 7666 1423 7710
<< via2 >>
rect 1386 7673 1416 7703
<< m2 >>
rect 1379 8066 1423 8110
<< m3 >>
rect 1379 8066 1423 8110
<< via2 >>
rect 1386 8073 1416 8103
<< m2 >>
rect 947 8066 991 8110
<< m3 >>
rect 947 8066 991 8110
<< via2 >>
rect 954 8073 984 8103
<< m2 >>
rect 947 7394 991 7438
<< m3 >>
rect 947 7394 991 7438
<< via2 >>
rect 954 7401 984 7431
<< m2 >>
rect 435 7394 479 7438
<< m3 >>
rect 435 7394 479 7438
<< via2 >>
rect 442 7401 472 7431
<< m2 >>
rect 435 7762 479 7806
<< m3 >>
rect 435 7762 479 7806
<< via2 >>
rect 442 7769 472 7799
<< m2 >>
rect 227 7762 271 7806
<< m3 >>
rect 227 7762 271 7806
<< via2 >>
rect 234 7769 264 7799
<< m2 >>
rect 227 7906 271 7950
<< m3 >>
rect 227 7906 271 7950
<< via2 >>
rect 234 7913 264 7943
<< m2 >>
rect 371 7906 415 7950
<< m3 >>
rect 371 7906 415 7950
<< via2 >>
rect 378 7913 408 7943
<< m2 >>
rect 371 7906 415 7950
<< m3 >>
rect 371 7906 415 7950
<< via2 >>
rect 378 7913 408 7943
<< m2 >>
rect 227 7906 271 7950
<< m3 >>
rect 227 7906 271 7950
<< via2 >>
rect 234 7913 264 7943
<< m2 >>
rect 227 7666 271 7710
<< m3 >>
rect 227 7666 271 7710
<< via2 >>
rect 234 7673 264 7703
<< m3 >>
rect 1243 6328 1273 7367
<< m2 >>
rect 1243 7337 1513 7367
<< m3 >>
rect 1483 7337 1513 8199
<< m2 >>
rect 1243 8169 1513 8199
<< m3 >>
rect 1243 8169 1273 8343
<< m3 >>
rect 1243 8313 1273 8343
<< m2 >>
rect 1099 8313 1273 8343
<< m3 >>
rect 1099 8313 1129 8519
<< m2 >>
rect 1099 8489 1273 8519
<< m3 >>
rect 1243 8489 1273 8743
<< m3 >>
rect 1243 8713 1273 8743
<< m2 >>
rect 1243 8713 1417 8743
<< m3 >>
rect 1387 8713 1417 9287
<< m2 >>
rect 1083 9257 1417 9287
<< m3 >>
rect 1083 9113 1113 9287
<< m2 >>
rect 811 9113 1113 9143
<< m3 >>
rect 811 8969 841 9143
<< m2 >>
rect 667 8969 841 8999
<< m3 >>
rect 667 8728 697 8999
<< m1 >>
rect 1205 8303 1315 8357
<< m2 >>
rect 1205 8303 1315 8357
<< via1 >>
rect 1212 8310 1308 8350
<< m1 >>
rect 1205 8303 1315 8357
<< m2 >>
rect 1205 8303 1315 8357
<< via1 >>
rect 1212 8310 1308 8350
<< m1 >>
rect 1205 8303 1315 8357
<< m2 >>
rect 1205 8303 1315 8357
<< via1 >>
rect 1212 8310 1308 8350
<< m1 >>
rect 1205 8703 1315 8757
<< m2 >>
rect 1205 8703 1315 8757
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 1205 8703 1315 8757
<< m2 >>
rect 1205 8703 1315 8757
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 1205 8703 1315 8757
<< m2 >>
rect 1205 8703 1315 8757
<< via1 >>
rect 1212 8710 1308 8750
<< m1 >>
rect 629 8703 739 8757
<< m2 >>
rect 629 8703 739 8757
<< via1 >>
rect 636 8710 732 8750
<< m1 >>
rect 1205 6303 1315 6357
<< m2 >>
rect 1205 6303 1315 6357
<< via1 >>
rect 1212 6310 1308 6350
<< m2 >>
rect 1236 7330 1280 7374
<< m3 >>
rect 1236 7330 1280 7374
<< via2 >>
rect 1243 7337 1273 7367
<< m2 >>
rect 1476 7330 1520 7374
<< m3 >>
rect 1476 7330 1520 7374
<< via2 >>
rect 1483 7337 1513 7367
<< m2 >>
rect 1476 8162 1520 8206
<< m3 >>
rect 1476 8162 1520 8206
<< via2 >>
rect 1483 8169 1513 8199
<< m2 >>
rect 1236 8162 1280 8206
<< m3 >>
rect 1236 8162 1280 8206
<< via2 >>
rect 1243 8169 1273 8199
<< m2 >>
rect 1236 8306 1280 8350
<< m3 >>
rect 1236 8306 1280 8350
<< via2 >>
rect 1243 8313 1273 8343
<< m2 >>
rect 1092 8306 1136 8350
<< m3 >>
rect 1092 8306 1136 8350
<< via2 >>
rect 1099 8313 1129 8343
<< m2 >>
rect 1092 8482 1136 8526
<< m3 >>
rect 1092 8482 1136 8526
<< via2 >>
rect 1099 8489 1129 8519
<< m2 >>
rect 1236 8482 1280 8526
<< m3 >>
rect 1236 8482 1280 8526
<< via2 >>
rect 1243 8489 1273 8519
<< m2 >>
rect 1236 8706 1280 8750
<< m3 >>
rect 1236 8706 1280 8750
<< via2 >>
rect 1243 8713 1273 8743
<< m2 >>
rect 1380 8706 1424 8750
<< m3 >>
rect 1380 8706 1424 8750
<< via2 >>
rect 1387 8713 1417 8743
<< m2 >>
rect 1380 9250 1424 9294
<< m3 >>
rect 1380 9250 1424 9294
<< via2 >>
rect 1387 9257 1417 9287
<< m2 >>
rect 1076 9250 1120 9294
<< m3 >>
rect 1076 9250 1120 9294
<< via2 >>
rect 1083 9257 1113 9287
<< m2 >>
rect 1076 9106 1120 9150
<< m3 >>
rect 1076 9106 1120 9150
<< via2 >>
rect 1083 9113 1113 9143
<< m2 >>
rect 804 9106 848 9150
<< m3 >>
rect 804 9106 848 9150
<< via2 >>
rect 811 9113 841 9143
<< m2 >>
rect 804 8962 848 9006
<< m3 >>
rect 804 8962 848 9006
<< via2 >>
rect 811 8969 841 8999
<< m2 >>
rect 660 8962 704 9006
<< m3 >>
rect 660 8962 704 9006
<< via2 >>
rect 667 8969 697 8999
<< m3 >>
rect 534 2018 564 2273
<< m2 >>
rect 534 2243 740 2273
<< m3 >>
rect 710 2243 740 2449
<< m2 >>
rect 710 2419 980 2449
<< m3 >>
rect 950 2419 980 2625
<< m2 >>
rect 950 2595 1140 2625
<< m3 >>
rect 1110 2595 1140 2785
<< m2 >>
rect 1110 2755 1284 2785
<< m3 >>
rect 1254 2755 1284 2977
<< m2 >>
rect 1254 2947 1460 2977
<< m3 >>
rect 1430 2947 1460 3265
<< m2 >>
rect 1430 3235 1700 3265
<< m3 >>
rect 1670 3235 1700 3409
<< m2 >>
rect 1670 3379 1860 3409
<< m3 >>
rect 1830 3379 1860 3553
<< m2 >>
rect 1830 3523 2020 3553
<< m3 >>
rect 1990 3523 2020 3857
<< m2 >>
rect 1990 3827 2277 3857
<< locali >>
rect 475 1953 633 2087
<< m1 >>
rect 475 1953 633 2087
<< viali >>
rect 482 1960 626 2080
<< locali >>
rect 2203 3773 2361 3907
<< m1 >>
rect 2203 3773 2361 3907
<< viali >>
rect 2210 3780 2354 3900
<< m2 >>
rect 527 2236 571 2280
<< m3 >>
rect 527 2236 571 2280
<< via2 >>
rect 534 2243 564 2273
<< m2 >>
rect 703 2236 747 2280
<< m3 >>
rect 703 2236 747 2280
<< via2 >>
rect 710 2243 740 2273
<< m2 >>
rect 703 2412 747 2456
<< m3 >>
rect 703 2412 747 2456
<< via2 >>
rect 710 2419 740 2449
<< m2 >>
rect 943 2412 987 2456
<< m3 >>
rect 943 2412 987 2456
<< via2 >>
rect 950 2419 980 2449
<< m2 >>
rect 943 2588 987 2632
<< m3 >>
rect 943 2588 987 2632
<< via2 >>
rect 950 2595 980 2625
<< m2 >>
rect 1103 2588 1147 2632
<< m3 >>
rect 1103 2588 1147 2632
<< via2 >>
rect 1110 2595 1140 2625
<< m2 >>
rect 1103 2748 1147 2792
<< m3 >>
rect 1103 2748 1147 2792
<< via2 >>
rect 1110 2755 1140 2785
<< m2 >>
rect 1247 2748 1291 2792
<< m3 >>
rect 1247 2748 1291 2792
<< via2 >>
rect 1254 2755 1284 2785
<< m2 >>
rect 1247 2940 1291 2984
<< m3 >>
rect 1247 2940 1291 2984
<< via2 >>
rect 1254 2947 1284 2977
<< m2 >>
rect 1423 2940 1467 2984
<< m3 >>
rect 1423 2940 1467 2984
<< via2 >>
rect 1430 2947 1460 2977
<< m2 >>
rect 1423 3228 1467 3272
<< m3 >>
rect 1423 3228 1467 3272
<< via2 >>
rect 1430 3235 1460 3265
<< m2 >>
rect 1663 3228 1707 3272
<< m3 >>
rect 1663 3228 1707 3272
<< via2 >>
rect 1670 3235 1700 3265
<< m2 >>
rect 1663 3372 1707 3416
<< m3 >>
rect 1663 3372 1707 3416
<< via2 >>
rect 1670 3379 1700 3409
<< m2 >>
rect 1823 3372 1867 3416
<< m3 >>
rect 1823 3372 1867 3416
<< via2 >>
rect 1830 3379 1860 3409
<< m2 >>
rect 1823 3516 1867 3560
<< m3 >>
rect 1823 3516 1867 3560
<< via2 >>
rect 1830 3523 1860 3553
<< m2 >>
rect 1983 3516 2027 3560
<< m3 >>
rect 1983 3516 2027 3560
<< via2 >>
rect 1990 3523 2020 3553
<< m2 >>
rect 1983 3820 2027 3864
<< m3 >>
rect 1983 3820 2027 3864
<< via2 >>
rect 1990 3827 2020 3857
<< m3 >>
rect 534 3840 564 4095
<< m2 >>
rect 534 4065 740 4095
<< m3 >>
rect 710 4065 740 4271
<< m2 >>
rect 710 4241 980 4271
<< m3 >>
rect 950 4241 980 4447
<< m2 >>
rect 950 4417 1140 4447
<< m3 >>
rect 1110 4417 1140 4607
<< m2 >>
rect 1110 4577 1284 4607
<< m3 >>
rect 1254 4577 1284 4799
<< m2 >>
rect 1254 4769 1460 4799
<< m3 >>
rect 1430 4769 1460 5087
<< m2 >>
rect 1430 5057 1700 5087
<< m3 >>
rect 1670 5057 1700 5231
<< m2 >>
rect 1670 5201 1860 5231
<< m3 >>
rect 1830 5201 1860 5375
<< m2 >>
rect 1830 5345 2020 5375
<< m3 >>
rect 1990 5345 2020 5695
<< m2 >>
rect 1990 5665 2277 5695
<< locali >>
rect 475 3773 633 3907
<< m1 >>
rect 475 3773 633 3907
<< viali >>
rect 482 3780 626 3900
<< locali >>
rect 2203 5623 2361 5757
<< m1 >>
rect 2203 5623 2361 5757
<< viali >>
rect 2210 5630 2354 5750
<< m2 >>
rect 527 4058 571 4102
<< m3 >>
rect 527 4058 571 4102
<< via2 >>
rect 534 4065 564 4095
<< m2 >>
rect 703 4058 747 4102
<< m3 >>
rect 703 4058 747 4102
<< via2 >>
rect 710 4065 740 4095
<< m2 >>
rect 703 4234 747 4278
<< m3 >>
rect 703 4234 747 4278
<< via2 >>
rect 710 4241 740 4271
<< m2 >>
rect 943 4234 987 4278
<< m3 >>
rect 943 4234 987 4278
<< via2 >>
rect 950 4241 980 4271
<< m2 >>
rect 943 4410 987 4454
<< m3 >>
rect 943 4410 987 4454
<< via2 >>
rect 950 4417 980 4447
<< m2 >>
rect 1103 4410 1147 4454
<< m3 >>
rect 1103 4410 1147 4454
<< via2 >>
rect 1110 4417 1140 4447
<< m2 >>
rect 1103 4570 1147 4614
<< m3 >>
rect 1103 4570 1147 4614
<< via2 >>
rect 1110 4577 1140 4607
<< m2 >>
rect 1247 4570 1291 4614
<< m3 >>
rect 1247 4570 1291 4614
<< via2 >>
rect 1254 4577 1284 4607
<< m2 >>
rect 1247 4762 1291 4806
<< m3 >>
rect 1247 4762 1291 4806
<< via2 >>
rect 1254 4769 1284 4799
<< m2 >>
rect 1423 4762 1467 4806
<< m3 >>
rect 1423 4762 1467 4806
<< via2 >>
rect 1430 4769 1460 4799
<< m2 >>
rect 1423 5050 1467 5094
<< m3 >>
rect 1423 5050 1467 5094
<< via2 >>
rect 1430 5057 1460 5087
<< m2 >>
rect 1663 5050 1707 5094
<< m3 >>
rect 1663 5050 1707 5094
<< via2 >>
rect 1670 5057 1700 5087
<< m2 >>
rect 1663 5194 1707 5238
<< m3 >>
rect 1663 5194 1707 5238
<< via2 >>
rect 1670 5201 1700 5231
<< m2 >>
rect 1823 5194 1867 5238
<< m3 >>
rect 1823 5194 1867 5238
<< via2 >>
rect 1830 5201 1860 5231
<< m2 >>
rect 1823 5338 1867 5382
<< m3 >>
rect 1823 5338 1867 5382
<< via2 >>
rect 1830 5345 1860 5375
<< m2 >>
rect 1983 5338 2027 5382
<< m3 >>
rect 1983 5338 2027 5382
<< via2 >>
rect 1990 5345 2020 5375
<< m2 >>
rect 1983 5658 2027 5702
<< m3 >>
rect 1983 5658 2027 5702
<< via2 >>
rect 1990 5665 2020 5695
<< m3 >>
rect 1244 8883 1274 9122
<< m2 >>
rect 1244 8883 1514 8913
<< m3 >>
rect 1484 8595 1514 8913
<< m2 >>
rect 1052 8595 1514 8625
<< m2 >>
rect 1244 9107 1562 9137
<< m3 >>
rect 1532 9107 1562 9281
<< m2 >>
rect 1532 9251 1706 9281
<< m3 >>
rect 1676 8995 1706 9281
<< m2 >>
rect 1052 8995 1706 9025
<< m3 >>
rect 1052 8995 1082 9025
<< m2 >>
rect 1052 8995 1610 9025
<< m3 >>
rect 1580 8995 1610 9505
<< m2 >>
rect 844 9475 1610 9505
<< m3 >>
rect 844 9315 874 9505
<< m2 >>
rect 508 9315 874 9345
<< m3 >>
rect 508 9139 538 9345
<< m2 >>
rect 284 9139 538 9169
<< m3 >>
rect 284 8995 314 9169
<< m2 >>
rect 284 8995 506 9025
<< m3 >>
rect 476 8595 506 9025
<< m2 >>
rect 140 8595 506 8625
<< m3 >>
rect 140 8355 170 8625
<< m2 >>
rect 140 8355 506 8385
<< m3 >>
rect 476 8195 506 8385
<< m3 >>
rect 476 8195 506 8225
<< m2 >>
rect 140 8195 506 8225
<< m3 >>
rect 140 7379 170 8225
<< m2 >>
rect 140 7379 314 7409
<< m3 >>
rect 284 7235 314 7409
<< m2 >>
rect 284 7235 1418 7265
<< m3 >>
rect 1388 7235 1418 7457
<< m2 >>
rect 1388 7427 1610 7457
<< m3 >>
rect 1580 7427 1610 7825
<< m2 >>
rect 1052 7795 1610 7825
<< m2 >>
rect 140 8195 506 8225
<< m3 >>
rect 140 7379 170 8225
<< m2 >>
rect 140 7379 314 7409
<< m3 >>
rect 284 7235 314 7409
<< m2 >>
rect 284 7235 1418 7265
<< m3 >>
rect 1388 7235 1418 7457
<< m2 >>
rect 1388 7427 1610 7457
<< m3 >>
rect 1580 7427 1610 7825
<< m2 >>
rect 1052 7795 1610 7825
<< m3 >>
rect 1052 7795 1082 7825
<< m2 >>
rect 1052 7795 1610 7825
<< m3 >>
rect 1580 7523 1610 7825
<< m2 >>
rect 1388 7523 1610 7553
<< m3 >>
rect 1388 7235 1418 7553
<< m2 >>
rect 1068 7235 1418 7265
<< m3 >>
rect 1068 7235 1098 7841
<< m2 >>
rect 844 7811 1098 7841
<< m3 >>
rect 844 7811 874 8225
<< m2 >>
rect 844 8195 1067 8225
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 7783 1123 7837
<< m2 >>
rect 1013 7783 1123 7837
<< via1 >>
rect 1020 7790 1116 7830
<< m1 >>
rect 1013 8183 1123 8237
<< m2 >>
rect 1013 8183 1123 8237
<< via1 >>
rect 1020 8190 1116 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 437 8183 547 8237
<< m2 >>
rect 437 8183 547 8237
<< via1 >>
rect 444 8190 540 8230
<< m1 >>
rect 1013 8583 1123 8637
<< m2 >>
rect 1013 8583 1123 8637
<< via1 >>
rect 1020 8590 1116 8630
<< m1 >>
rect 437 8583 547 8637
<< m2 >>
rect 437 8583 547 8637
<< via1 >>
rect 444 8590 540 8630
<< m1 >>
rect 437 8583 547 8637
<< m2 >>
rect 437 8583 547 8637
<< via1 >>
rect 444 8590 540 8630
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 1013 8983 1123 9037
<< m2 >>
rect 1013 8983 1123 9037
<< via1 >>
rect 1020 8990 1116 9030
<< m1 >>
rect 437 8983 547 9037
<< m2 >>
rect 437 8983 547 9037
<< via1 >>
rect 444 8990 540 9030
<< m1 >>
rect 437 8983 547 9037
<< m2 >>
rect 437 8983 547 9037
<< via1 >>
rect 444 8990 540 9030
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m1 >>
rect 1205 9103 1315 9157
<< m2 >>
rect 1205 9103 1315 9157
<< via1 >>
rect 1212 9110 1308 9150
<< m2 >>
rect 1237 8876 1281 8920
<< m3 >>
rect 1237 8876 1281 8920
<< via2 >>
rect 1244 8883 1274 8913
<< m2 >>
rect 1477 8876 1521 8920
<< m3 >>
rect 1477 8876 1521 8920
<< via2 >>
rect 1484 8883 1514 8913
<< m2 >>
rect 1477 8588 1521 8632
<< m3 >>
rect 1477 8588 1521 8632
<< via2 >>
rect 1484 8595 1514 8625
<< m2 >>
rect 1525 9100 1569 9144
<< m3 >>
rect 1525 9100 1569 9144
<< via2 >>
rect 1532 9107 1562 9137
<< m2 >>
rect 1525 9244 1569 9288
<< m3 >>
rect 1525 9244 1569 9288
<< via2 >>
rect 1532 9251 1562 9281
<< m2 >>
rect 1669 9244 1713 9288
<< m3 >>
rect 1669 9244 1713 9288
<< via2 >>
rect 1676 9251 1706 9281
<< m2 >>
rect 1669 8988 1713 9032
<< m3 >>
rect 1669 8988 1713 9032
<< via2 >>
rect 1676 8995 1706 9025
<< m2 >>
rect 1045 8988 1089 9032
<< m3 >>
rect 1045 8988 1089 9032
<< via2 >>
rect 1052 8995 1082 9025
<< m2 >>
rect 1045 8988 1089 9032
<< m3 >>
rect 1045 8988 1089 9032
<< via2 >>
rect 1052 8995 1082 9025
<< m2 >>
rect 1573 8988 1617 9032
<< m3 >>
rect 1573 8988 1617 9032
<< via2 >>
rect 1580 8995 1610 9025
<< m2 >>
rect 1573 9468 1617 9512
<< m3 >>
rect 1573 9468 1617 9512
<< via2 >>
rect 1580 9475 1610 9505
<< m2 >>
rect 837 9468 881 9512
<< m3 >>
rect 837 9468 881 9512
<< via2 >>
rect 844 9475 874 9505
<< m2 >>
rect 837 9308 881 9352
<< m3 >>
rect 837 9308 881 9352
<< via2 >>
rect 844 9315 874 9345
<< m2 >>
rect 501 9308 545 9352
<< m3 >>
rect 501 9308 545 9352
<< via2 >>
rect 508 9315 538 9345
<< m2 >>
rect 501 9132 545 9176
<< m3 >>
rect 501 9132 545 9176
<< via2 >>
rect 508 9139 538 9169
<< m2 >>
rect 277 9132 321 9176
<< m3 >>
rect 277 9132 321 9176
<< via2 >>
rect 284 9139 314 9169
<< m2 >>
rect 277 8988 321 9032
<< m3 >>
rect 277 8988 321 9032
<< via2 >>
rect 284 8995 314 9025
<< m2 >>
rect 469 8988 513 9032
<< m3 >>
rect 469 8988 513 9032
<< via2 >>
rect 476 8995 506 9025
<< m2 >>
rect 469 8588 513 8632
<< m3 >>
rect 469 8588 513 8632
<< via2 >>
rect 476 8595 506 8625
<< m2 >>
rect 133 8588 177 8632
<< m3 >>
rect 133 8588 177 8632
<< via2 >>
rect 140 8595 170 8625
<< m2 >>
rect 133 8348 177 8392
<< m3 >>
rect 133 8348 177 8392
<< via2 >>
rect 140 8355 170 8385
<< m2 >>
rect 469 8348 513 8392
<< m3 >>
rect 469 8348 513 8392
<< via2 >>
rect 476 8355 506 8385
<< m2 >>
rect 469 8188 513 8232
<< m3 >>
rect 469 8188 513 8232
<< via2 >>
rect 476 8195 506 8225
<< m2 >>
rect 133 8188 177 8232
<< m3 >>
rect 133 8188 177 8232
<< via2 >>
rect 140 8195 170 8225
<< m2 >>
rect 133 7372 177 7416
<< m3 >>
rect 133 7372 177 7416
<< via2 >>
rect 140 7379 170 7409
<< m2 >>
rect 277 7372 321 7416
<< m3 >>
rect 277 7372 321 7416
<< via2 >>
rect 284 7379 314 7409
<< m2 >>
rect 277 7228 321 7272
<< m3 >>
rect 277 7228 321 7272
<< via2 >>
rect 284 7235 314 7265
<< m2 >>
rect 1381 7228 1425 7272
<< m3 >>
rect 1381 7228 1425 7272
<< via2 >>
rect 1388 7235 1418 7265
<< m2 >>
rect 1381 7420 1425 7464
<< m3 >>
rect 1381 7420 1425 7464
<< via2 >>
rect 1388 7427 1418 7457
<< m2 >>
rect 1573 7420 1617 7464
<< m3 >>
rect 1573 7420 1617 7464
<< via2 >>
rect 1580 7427 1610 7457
<< m2 >>
rect 1573 7788 1617 7832
<< m3 >>
rect 1573 7788 1617 7832
<< via2 >>
rect 1580 7795 1610 7825
<< m2 >>
rect 133 8188 177 8232
<< m3 >>
rect 133 8188 177 8232
<< via2 >>
rect 140 8195 170 8225
<< m2 >>
rect 133 7372 177 7416
<< m3 >>
rect 133 7372 177 7416
<< via2 >>
rect 140 7379 170 7409
<< m2 >>
rect 277 7372 321 7416
<< m3 >>
rect 277 7372 321 7416
<< via2 >>
rect 284 7379 314 7409
<< m2 >>
rect 277 7228 321 7272
<< m3 >>
rect 277 7228 321 7272
<< via2 >>
rect 284 7235 314 7265
<< m2 >>
rect 1381 7228 1425 7272
<< m3 >>
rect 1381 7228 1425 7272
<< via2 >>
rect 1388 7235 1418 7265
<< m2 >>
rect 1381 7420 1425 7464
<< m3 >>
rect 1381 7420 1425 7464
<< via2 >>
rect 1388 7427 1418 7457
<< m2 >>
rect 1573 7420 1617 7464
<< m3 >>
rect 1573 7420 1617 7464
<< via2 >>
rect 1580 7427 1610 7457
<< m2 >>
rect 1573 7788 1617 7832
<< m3 >>
rect 1573 7788 1617 7832
<< via2 >>
rect 1580 7795 1610 7825
<< m2 >>
rect 1045 7788 1089 7832
<< m3 >>
rect 1045 7788 1089 7832
<< via2 >>
rect 1052 7795 1082 7825
<< m2 >>
rect 1045 7788 1089 7832
<< m3 >>
rect 1045 7788 1089 7832
<< via2 >>
rect 1052 7795 1082 7825
<< m2 >>
rect 1573 7788 1617 7832
<< m3 >>
rect 1573 7788 1617 7832
<< via2 >>
rect 1580 7795 1610 7825
<< m2 >>
rect 1573 7516 1617 7560
<< m3 >>
rect 1573 7516 1617 7560
<< via2 >>
rect 1580 7523 1610 7553
<< m2 >>
rect 1381 7516 1425 7560
<< m3 >>
rect 1381 7516 1425 7560
<< via2 >>
rect 1388 7523 1418 7553
<< m2 >>
rect 1381 7228 1425 7272
<< m3 >>
rect 1381 7228 1425 7272
<< via2 >>
rect 1388 7235 1418 7265
<< m2 >>
rect 1061 7228 1105 7272
<< m3 >>
rect 1061 7228 1105 7272
<< via2 >>
rect 1068 7235 1098 7265
<< m2 >>
rect 1061 7804 1105 7848
<< m3 >>
rect 1061 7804 1105 7848
<< via2 >>
rect 1068 7811 1098 7841
<< m2 >>
rect 837 7804 881 7848
<< m3 >>
rect 837 7804 881 7848
<< via2 >>
rect 844 7811 874 7841
<< m2 >>
rect 837 8188 881 8232
<< m3 >>
rect 837 8188 881 8232
<< via2 >>
rect 844 8195 874 8225
<< locali >>
rect 100 9840 2736 9890
<< locali >>
rect 100 100 2736 150
<< m1 >>
rect 100 150 150 9840
<< m1 >>
rect 2686 150 2736 9840
<< locali >>
rect 93 9833 157 9897
<< m1 >>
rect 93 9833 157 9897
<< viali >>
rect 100 9840 150 9890
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 2679 9833 2743 9897
<< m1 >>
rect 2679 9833 2743 9897
<< viali >>
rect 2686 9840 2736 9890
<< locali >>
rect 2679 93 2743 157
<< m1 >>
rect 2679 93 2743 157
<< viali >>
rect 2686 100 2736 150
<< locali >>
rect 0 9940 2836 9990
<< locali >>
rect 0 0 2836 50
<< m1 >>
rect 0 50 50 9940
<< m1 >>
rect 2786 50 2836 9940
<< locali >>
rect -7 9933 57 9997
<< m1 >>
rect -7 9933 57 9997
<< viali >>
rect 0 9940 50 9990
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 2779 9933 2843 9997
<< m1 >>
rect 2779 9933 2843 9997
<< viali >>
rect 2786 9940 2836 9990
<< locali >>
rect 2779 -7 2843 57
<< m1 >>
rect 2779 -7 2843 57
<< viali >>
rect 2786 0 2836 50
<< locali >>
rect 828 9390 1116 9430
<< locali >>
rect 252 9390 540 9430
<< locali >>
rect 636 9270 796 9310
<< locali >>
rect 252 6590 540 6630
<< locali >>
rect 636 6470 796 6510
<< locali >>
rect 828 6590 1116 6630
<< locali >>
rect 100 7322 2736 7418
<< locali >>
rect 93 7315 157 7425
<< m1 >>
rect 93 7315 157 7425
<< viali >>
rect 100 7322 150 7418
<< locali >>
rect 2679 7315 2743 7425
<< m1 >>
rect 2679 7315 2743 7425
<< viali >>
rect 2686 7322 2736 7418
<< locali >>
rect 100 9562 2736 9658
<< locali >>
rect 93 9555 157 9665
<< m1 >>
rect 93 9555 157 9665
<< viali >>
rect 100 9562 150 9658
<< locali >>
rect 2679 9555 2743 9665
<< m1 >>
rect 2679 9555 2743 9665
<< viali >>
rect 2686 9562 2736 9658
<< locali >>
rect 0 6762 2836 6858
<< locali >>
rect -7 6755 57 6865
<< m1 >>
rect -7 6755 57 6865
<< viali >>
rect 0 6762 50 6858
<< locali >>
rect 2779 6755 2843 6865
<< m1 >>
rect 2779 6755 2843 6865
<< viali >>
rect 2786 6762 2836 6858
<< locali >>
rect 0 6122 2836 6218
<< locali >>
rect -7 6115 57 6225
<< m1 >>
rect -7 6115 57 6225
<< viali >>
rect 0 6122 50 6218
<< locali >>
rect 2779 6115 2843 6225
<< m1 >>
rect 2779 6115 2843 6225
<< viali >>
rect 2786 6122 2836 6218
<< locali >>
rect 308 5630 626 5750
<< locali >>
rect 0 2164 2836 2220
<< locali >>
rect -7 2157 57 2227
<< m1 >>
rect -7 2157 57 2227
<< viali >>
rect 0 2164 50 2220
<< locali >>
rect 2779 2157 2843 2227
<< m1 >>
rect 2779 2157 2843 2227
<< viali >>
rect 2786 2164 2836 2220
<< locali >>
rect 0 500 2836 556
<< locali >>
rect -7 493 57 563
<< m1 >>
rect -7 493 57 563
<< viali >>
rect 0 500 50 556
<< locali >>
rect 2779 493 2843 563
<< m1 >>
rect 2779 493 2843 563
<< viali >>
rect 2786 500 2836 556
<< locali >>
rect 0 3984 2836 4040
<< locali >>
rect -7 3977 57 4047
<< m1 >>
rect -7 3977 57 4047
<< viali >>
rect 0 3984 50 4040
<< locali >>
rect 2779 3977 2843 4047
<< m1 >>
rect 2779 3977 2843 4047
<< viali >>
rect 2786 3984 2836 4040
<< locali >>
rect 0 2320 2836 2376
<< locali >>
rect -7 2313 57 2383
<< m1 >>
rect -7 2313 57 2383
<< viali >>
rect 0 2320 50 2376
<< locali >>
rect 2779 2313 2843 2383
<< m1 >>
rect 2779 2313 2843 2383
<< viali >>
rect 2786 2320 2836 2376
<< locali >>
rect 0 5834 2836 5890
<< locali >>
rect -7 5827 57 5897
<< m1 >>
rect -7 5827 57 5897
<< viali >>
rect 0 5834 50 5890
<< locali >>
rect 2779 5827 2843 5897
<< m1 >>
rect 2779 5827 2843 5897
<< viali >>
rect 2786 5834 2836 5890
<< locali >>
rect 0 4170 2836 4226
<< locali >>
rect -7 4163 57 4233
<< m1 >>
rect -7 4163 57 4233
<< viali >>
rect 0 4170 50 4226
<< locali >>
rect 2779 4163 2843 4233
<< m1 >>
rect 2779 4163 2843 4233
<< viali >>
rect 2786 4170 2836 4226
<< locali >>
rect -100 10040 2936 10090
<< locali >>
rect -100 -100 2936 -50
<< m1 >>
rect -100 -50 -50 10040
<< m1 >>
rect 2886 -50 2936 10040
<< locali >>
rect -107 10033 -43 10097
<< m1 >>
rect -107 10033 -43 10097
<< viali >>
rect -100 10040 -50 10090
<< locali >>
rect -107 -107 -43 -43
<< m1 >>
rect -107 -107 -43 -43
<< viali >>
rect -100 -100 -50 -50
<< locali >>
rect 2879 10033 2943 10097
<< m1 >>
rect 2879 10033 2943 10097
<< viali >>
rect 2886 10040 2936 10090
<< locali >>
rect 2879 -107 2943 -43
<< m1 >>
rect 2879 -107 2943 -43
<< viali >>
rect 2886 -100 2936 -50
<< locali >>
rect -200 10140 3036 10190
<< locali >>
rect -200 -200 3036 -150
<< m1 >>
rect -200 -150 -150 10140
<< m1 >>
rect 2986 -150 3036 10140
<< locali >>
rect -207 10133 -143 10197
<< m1 >>
rect -207 10133 -143 10197
<< viali >>
rect -200 10140 -150 10190
<< locali >>
rect -207 -207 -143 -143
<< m1 >>
rect -207 -207 -143 -143
<< viali >>
rect -200 -200 -150 -150
<< locali >>
rect 2979 10133 3043 10197
<< m1 >>
rect 2979 10133 3043 10197
<< viali >>
rect 2986 10140 3036 10190
<< locali >>
rect 2979 -207 3043 -143
<< m1 >>
rect 2979 -207 3043 -143
<< viali >>
rect 2986 -200 3036 -150
<< labels >>
flabel m2 s 969 7673 1416 7703 0 FreeSans 400 0 0 0 INP
port 1 nsew signal bidirectional
flabel m2 s 234 8473 393 8503 0 FreeSans 400 0 0 0 INN
port 2 nsew signal bidirectional
flabel locali s 100 9840 2736 9890 0 FreeSans 400 0 0 0 VDD
port 3 nsew signal bidirectional
flabel locali s 0 9940 2836 9990 0 FreeSans 400 0 0 0 VSS
port 4 nsew signal bidirectional
flabel m3 s 1243 6328 1273 7367 0 FreeSans 400 0 0 0 OUT
port 5 nsew signal bidirectional
flabel locali s -100 10040 2936 10090 0 FreeSans 400 0 0 0 VDD
port 48 nsew signal bidirectional
flabel locali s -200 10140 3036 10190 0 FreeSans 400 0 0 0 VSS
port 49 nsew signal bidirectional
<< properties >>
<< end >>